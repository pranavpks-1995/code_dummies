package Code_Generator;
	module program (Empty);
	endmodule
endpackage