���)ޛ}(�Qp�w�;����ێ���v�u�c��O��_Ɇ�t����;=x�]P2���Z������RL���؝%ń<D#�s�+u�Nt�a���c{&����Rn=��d��4�4Q"r�X���A�y۶/n��/��KH?霨��bb�;�8�"��1�LSd��׊��Mm� �ZhC�r���̂6�pX��a��?໘����f�E0�0�&��8�إ��ۑ�\`̃�T���b���~��;4�t�o��CS�w�׻9�C�Ds���Uz����.�q��R�|���BV2����5��J@OO��`�.-5�Q�ڪT�b{wo�^���C0M|�e�l�R�D���|���iw+�<;)�.�`���F4��2���@���e��@=�kY��s�<�tM�����حe�4�]�����MhI8���+����;��\]�92�I�n�y+��-��'`���9p�<*gp��D����]�<�A�-����� $�KOJ>�L� �[�'�gD��c#P�������[�����`	}��8[ =��k�%(�2=�����}wIu>ໄ'�KP������MЏ�?�ٞq*�5f��@��t�7�&L���Q�Z�E�_O9wƑ����㭊`������*8��Ͻ����%Ħo�� ����Q�Z��9�Ff5��VQ�~W�R�,�$��כ#<�ݍ�}��3ۛik�0j&��@D����>l��\C��@���fX��"���!�<Uiw�3vR�'��
��<Nd@�H�$�?��<����I@�\�E����I2��G �a��K���I�G��}_Ԩ�P�?��L���"��m�*��wC\���>n�.������L�Qxb�!��Y����x��]=�^�@��z�w>1�"��������nv����{Y鎏�3B .\���e&��!t����~��0����#��{�i�ߒ�nq��*z����]�vN����h�^j��Ox��pw��[iv�3�%��L�ǝ��%Ӓⲗ��������\T����YL�s�O������B1.�0*��,Z
7Yb�%��i��o��@ׇb�&H����r}�����T��X-��(�j|:l���B�(�ٞư��E���;
ll%T�h4����8�r��;a���.-]�ܶ6���G�,�8�Рâ:�{V�{���
������h�A�:��@@a\#r�n��i���)#���%��=u���_)86���h��?B |��DN�o���'0�e�.O����_E҈5�"�vw8:0mÇ��p$�����D��(�iKtb���G�o	mV,4H�J%��o�:�������f�w{��4�I�c�Q���ǳ�*a��hˡ����)b���<0���q#��ށ�g�Q
Nk�P���pi	ϵZ}#��.25zB�X�(���;�3ʽѼϞ�e���f��eU
�tZ����IK�j�}��n�AK���r�6�kW&�>�ۺ`2X������
2gE�����mF����3XcM-���*ٺ����-;��X��n�I�{�B��jD�����=0���������/\�bt�;�B?����s�<r�8`��=�	��FH�{X$6���V��Վ��,�	ԕ�Jm�����-2��WO5q�:�$'� �'ܨ��E1q�xD�ogr��S��֚���4J��2�	o� Q	��&o
<Q"x.�����zr|����RK$Y��6��V�;���v�3��>Jt9M��@&��!ÊMA5�W&x���V+B�"�5��r��Wf�!-Ca1[B����r/-�X�
H�x+XȦ��G��.�������B9'�Vib��;�vO�#�(��|�� {?&�~�mTx����z����ȬD%D����{��Y4�4���0���x ���֖ͤ9D�4l����IKB�P�j���gPj� �9&ۯC�}r�>M�3Wh�!U�V�%�õ����'V�mv`�KR��p]XW	��J�3;�H�k��sK����[ �s����+���b�t]
�}��ǔ�>e�C�q�w|$�R��!�辪��A=�@-MW>?ځT%I>�KY���i�M�����+ޏl���X��k���EY��-'��$'�8#�Pf'r֯�l��x������%US�Օ��qj_���w�W��r��qY���
��1�?��v�3�
��I�������2
�Զ�^����p���W<l���@B����X�D`����w��^��j������Y��A]�M�u������(�a��C��[ E�Fԑ��7=x����Xp�0��C'������ˤ&!���s<I�N�X�]��g�le�#�3�+�@nDd.���Tt��$[�zi��?��4���g��'b�RS��$!����:Q�����Y��{ώ�_8İ��]�2��x�v�Dbwݣ�4L��P^ ���1�H�u��wf�3�,�Pi�Z$�,TZ�U^u;����'�`^3~�)�5��)k�-���rYarF�Zg�~�G}צ���fl�)�Tf����|��:�*�Fc*�^ێʹ��4�	��>��9R��"]𒜖��;V��8�,J=�����GDԒ ��F�� �8S�r�� 	W�0h����N��