B��@�q����)<"�Vr���Ff��F� �1
��g}�ߎ!�g(V9n�f������n  !K�GRbT]4��7Q�2X�xf,����z�V#0�Jl�L	�O(�S�F�Xl�.ܕ�Ɖ��{���&�2U���(X��!`m�B��(�0vicR�a7J��-�xP��㐅C9/�-��5d�hp-wW��pb�R6%����y9E]��"L�A"�G�a�>i��#� O�hC���YN�@���.}F�^Ax 
�⹱�u����<�۵�[�4�UR�H�͖��    8!y������8�@�T �����Uy����4��'}OD��L�|�mR��8�]�Y"A��\T.�[K/�eӉ�&m���-��H3]�J��0ˌ��F��T:S#�,P��*��0�5�=�>\�J�@��)�"" E�D�M��^��r����$���YhV��[��U�c-� �     �!��IP�0�)2k4�@ C�m��D�2�X�t�"���f��%�k{�sMM�vW$lѥ -��[md��ޅ� h* ����Z��?wA�	̥�Gv��V��| Q�)ʌ�Gޢ.����h9��� ���ϐX��@ ���>�W�E�i�����e��ɖ��    �!��0�ga!"a�$h��J�p�O~AA�-c�����@��b�ORtx���؎�� �����O�.�V�u��� (�X��R���8jyٌs�Qy���$�;�>�1�.���B�gy%H���RY��۞P�P��'g�W�$��zFn��'n�> `    !)��0��P� h
�wi�
�Bv��e�^�l�U;�[��Z# �gr�
�= ?½]���2�����eS��\]�k]J�I��}eM���$�׵��c��`3aJðrF����o5��,�� Ȥ"!�`P`rr�Gx����$��+cf `    !K�GCNi�(��aWR
�*����@UZ�