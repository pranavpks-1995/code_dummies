�EJ��H�^`Ȱ��4�h���m�.�f���%�г��SCNʓ�fb�q���Ac��Mc|�_������}<xE����F� 6P1��x��*r: �*5�J�%I\8`��UoZҾBB;��G�����Rܖ�8�r��+;$�[����`zg�>��6�k�t���^c:	��U\a��N�O�����re��(�K2J�Z�[m^Iӳ�0�3�D;>��`��J�͹
�}8�-���E�܂�_�1L󟷈��DK��V
�ܦ ��5�-b8�����W���c��ܚE��x˭p[G��!e�9i��F����"qٙE/��/�~m���p.̍ n	#�4F]6���i�uh�?�2�����5z^�P��\�p�j�܅�vJ��~��%��a8
�.0�P�K�����W���/�Zj��7�ʸ�U�o��/��zH0���[Y����$�n9N��P%vh�3���Ԋ�<�;}� ����DՈS�:�����LZU��:�٢����ýE�s��4��+ ��p�1���jt�0����6_�]" P��Lɟ��$m����c,
��:+Kܦ*w��%&FoSI<����%�rZ�e~���X������w�E�t�����)2���z��1�P�\��������Sk8�W-��yw�V+'�Jn����m�gM ��|��ٵ��Ғ�@���U4fbbj�WZUc���fF�L���&D���c�K�yHX�� �O���$�f�e��M�q�r:�E� �ݜC��膭��ԗ�3��{�I3�YP���G�Z�RE[��F�aج#Y<].d��F`��G���i,�Zu�֒��cLh~��������H"�4r��V^�tK�7� ��f�X��M��7E1mJ<�0�I���DL�و"�C�M�
]�5�R�1�p�|�!	0�ےہ��_	�o�)�j�Z�����h�,�3g��yT�g�m'd�+h���	����cW���rHjQJ�|�ϥ�w;��~�st���'QX��>�4�af)��o�����bdW3�"1X=��������E�l���H���c͹�����_�u$P�:7�&ǵF0ݧ�;C��^��nyDYN8��Ny�Q�N�H�0<3�+�8]��'�n���S��m��i0̮Ұ�}��n�c^�,�l2� ��U47P����r��KPs����=|���o�C�C��Aw>��f[����A���'��yws���b���'���O��D����0p��g�1�.V�[����n�'�fT\0��m��ڴ�Bd�J���Pb�\bѢ���"E��۬��o��o�f�D,���k�r�;[Yݨ)�uWԯ���\�Y�'ï5���<�߀)�T0�Ij��B/�ê��kHW�A���c�K�=�J�+Di���*�@�C
������3�"4��;��]X��M=5T�����ϼ	� A�&Al�C���F����^������8 �����ե%y��D���l@��`�p3X!WT"��<��������$b��޽aC��9C��'w���MIs�zݮ��}'����O �<37�y����> 
^w�^v�W���G`N��-�R�ZפW�V��>�P����*n���9L��At�`��;�S"������l��P昪)K�2Wu�0 Ax����wۛ�[kM����k�}�@�lE���Ps���)4)_r�jn��[�k�����W�Nt��jY�ny���y���a���IM�vU]��A���n�&����`��M������֢���v���AsI��,�T���� B�������^��gs�������4�.��k	e\K�8KAn@�κ٭p]�W�M��3�p%���'��H���u�nFi[�1�ȩ��:x�5h��+��Hxﱬ�\��J��>��9a����9&�5�ZGU��ݎ�:���sUo�����'%6��BID5��PL�a(������Yzc����k�`�m<�d��M�S��}��'$�F�R��(�5����r��靶Jx���+wR*6?�����~R��wR%�n�"��|�K���i�����*��4�;'u��y�A�)$�8殦�����\�D⟏"Ri�̯����O;:8�i=����$��y5U�z4}"w�ψ�~0�B���u����fn���w��&���,����7�.�#�����qX�T���<�#���h�N3Im&�gd�mo���Wd �:�<���o�Lb^:�`Vr��[薡R��X;BK��z���WQ�[����N��+(����H�6']��'#d� �i֚Y�`���N�ۿ�����%��E�Kƛ֡r���ԩ��M�����?2=�2]�;�(��vܾ/uz�SG��}hEt$Oh�wR�ɍ��S�tGa�;��4[7�$�4�oV"��]��,�v��1��p�nm�r���/�C�tq��[���+��PȤ�|��㑗d��p�%ǰ6ˢ�4���H0�
�i��|fU��lS%Oͣ�kETG5<���<��	
���7�^���5�����<�)(h�h��$ǽ�0����?y��ǰ�y��$}v�ӗ�@�oE�Kq��1;����5qGOG�,��H����0�]_n�W����n���PB�!�5S�P���ؙ�D`��s���1�F$ZD����r����}����AG	!�%/�s��s��n:J{奌��1g�2<pP@������Hx��I}���p�D	�#�����X��*��p��F0���P��.�V�����{���]Nn�%�!Vz�5O�&/����B��K�U�)Ά����a��M��N��):�)�5��cr�Fu�|�p,Y�5p*��@s�\׌>��C�=,��o��H�犦�v�����a� ���&���YG�����ǹ�3%k�	���U���h���r��Q��J�_0b�=qf�)c�أ>�kS����7.w������$��k�����������.����9���L��Q��O��6�J͝���2����,V�Qk��S�|I��N��z��E���Q����&P1-���ɵ���lV±O�J3������&��e�[�����W����G�#������q��K��F����{���]p���Ce;�@|7��mm���n����g�,�߬\-ܻ�#�5���y#)���`����@m&�Q���"�V��V���!�W�V��Nj�}�(��|�ZN*Ai�@,8�����O�me��AhK�	��!}9`Q�������GO@�C�:)P�~D&Co�U�-S��B�^�X ѯ�aX�/�~�\[�i�����B|D�*��0v�k�z�)�|'��Q6e��262/�c��^�]Ux=��ƹ�x�]��3���Jk�����V[�J�с�P�2�X��4���h�w�KG����R�X�FA^0�:"����Ekb������"&�
X=��LFE�if"��������7no�a��3e�f\m@�ڐ���q������\
�m��;�TzEO�����N(�t�r��ߑ7:|%�1J���c��0R0]��hg���ͫ��l���5�t�\��O(��/l��5Z1+���p��4��T�@#����8��]���7_��y�me��V/^�4��"4{]��4�����"����RhN��:�sѕP.��h�`�"c"�a+k�LX!�w���8�M��4ID�kR}}@@��Kk���ҡj�0�����5�"�'JP(��JA��ZEWi�)_��j?x�����%7Hx�,�x�������Ȗ� �0�8����� x�ƞ�p�1w��S{���;�j����m��7�*����fe5����G~���g<��!x8|5��]���I����M?􊹏v�����B�㺏�c��	�:���.�ԇ��zqN�l�77_�'Z�p�B�KT�h��O����`�� ��x�+kmo�sm8GA<�&�z<0�]&<n��oc�[�XCe;v{9-K]�qk��1R����L�)�q��a)6OȞ�wa�ѻ��(������q�~lx,h�'�����)"�~�4��ږ�˽0IuQN�02�v�c���2���/U�Ħன	'�ʋƏv������>��[}8`�A���v>S䐂�Ơr*�J��ˋg?��-P�-w�ȥ���"&6!� ����"�z\��y��Ւ��42F�2@���7���x�5���~'��V�ew(�m`�k(K/��en��1E��Q]8H
i*�Z5�l���uQ�\�~�C"��w��(a83X���a8V��3�����0׵����Q�@����?��י�M�e���mc�}\��C�����&�(�v�,3��씯�
�y�k����V2
���x�ÍUI4b���#�TW"}8�:���2�a ���Z�jj��6p ���]R(��w���#��*5Я'FYF^^�8�j��<L�"8"�W�����[��=&��G�
=8ņR�}փ���������}��3czȬ���G�����g�`�Ô"8��uzi���V��]v���6�������a�9s鼠8(^l��3�~".������H8Oy�����䒤�5�qD ���R�&�h��؜�_�V�x���ݭ�R�C�l-v���7{��u�Nn��k2�}�эS|Sé�uR�f#��51��|��+W������(N��!���x���W���87�8�U4�.�� ��'|Y�n,*2�x��aq��V��&��yPM
!Ŋ)�ͼ��6�������C��X��G��K����a�ql��fΜh���0D�n��.,���J����x�d2&����2��^h���`ּH��f���w[����
U�Q��o���SvO_]���j�F9�ĺ��ީ�F�W-jXL1��Q�����JA�m��Ž��c��9� E ��)X���թ�ðK�-N[U\��G��9���O=Rr�C.��F���C�`�e��E�(pD�ɲ5V��u�DO��a�{0�S��I�c�O�h�2O�)6�c��w�
�ى_�_f'���m� ��r���l��?W}Dr ���b�%�T��b��He�_�`�>آ�*(�bu9�5��9Cr�t`n;fς�%�w�H��S �`i���o��ny<B���ľ�(�= J�ˏ��C2�V�3K�y�
D��ɏ���#!�O-����U+Кqlm�K�	
��eD�K�b3B�.�,|~~��R��9=R�v�|�+ϾK#_g:�_Wȓe��+�K�J�)+.�_#��*.�W]:9�z�E#��	�]{�B|��=c5�@�d�,I�Eg����е,���?J�Sր�%�} ]�v[{�A�:��-G�9d�����q�=s�Kr�����a��Ki١	I�#
دk�V�.�g��E�̖jJ�8m=8��5�T�s��X锼���gz����<�0P	S	��RxP��C�F5�8�Rr�s�i��9�#N���(8�ߓ9��Rep��1����jM��բ������uL����T�C�`?�I�釔,j%I�"����_��o�Iѓg����y�3\��C��o��PS05���7촟�o��b��G�ߴ�J@:�:�H�P���↹5�֘_vmS.�+�n�xum����X3�A���I����М�����e�%����uKY��M^*��v��\-h�8���6l��-����ڐ��+��k�6�J�V�f'��I���y�7x��1�{D�:ܗ�A��e�����q[�ܗp���q��	:��f�s0�I�#z��.�ɥ�������`؛�e��l�)Q C��6�W���/�A��`�.�.LV̱u��P#n��^���L�VlthrY$3��q�m�b�ܔ�[".Ɓ����|��5t�^���c��:p���5���Zq�>�ؤ6��Z�J\BA�5���Σw�����(�&��+���B�Yio�W����W���C�E�ae;ҟTÕ��ɎX ��M-��'I�|����O}ԃ��0�٘�<b�cwnC�mSX��yq���!��6�9ea��QlG�9�7�\�oHV�������}��2����ߟ2lˁ�z���j�X}e�qo��ƍ�.Ita�MU`�
�'�P������9����hoF�ds?PM�M)u˿�c�:�p|��M�+�L��ECP�U����16W�#�?��O�o_�d
�&S8��ov\=2=��˸�Pu3�,�g�vg�&��g?�5�s)�V(R_�SQ,�2�N"2 _W=