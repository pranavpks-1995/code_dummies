`��؎E�aF�i��jq�J2D����i�[���1j� 0����3s�i�- ��O�5O����R��y�N����[��wf\�q������|I��5���Ɣz-}��r���Ż��zH�?l"ҿV핇5����X�э�x_5I�J'	$���\1�������r��� ��s^)����p��K���$��%@�v���B�d��S6|��c�\���_Fc�i.`B/:c�w%~�ô��R1�*�W)���æ�g>>�Sˑ�ez��U���d��D�A�G�I���ƿ��p/�z�0�s��zq%�Ɨ:wK����[dP���°�أk�5$eC��z�X� ��7H�8m�ē>�Kv��*k�� ]�%f-���f&�8���9��"y?�w�����!���7v��4:$�� pOq4S�-�N�l2��
|��x,�̓�[�輳=�°lי$622�V�}S�o#Eׂ���Uvh�!<�SĢ-\���Z��-c`,������S�g"��E�����S��*��GCY?[��c1�ݪ�I�2�꠺^���V21����8��$v���2�A%��ܡ��s�I�wR�i35�iR���F���o�κ�7�GB�*ț�����DN�G$s�;,����g�ó��n�`���nI�P�Gc��:�A���=�z0/-FG��>9�Ov�֏���c��b2@���
�G_O=h.�u�ːnٵ�����I'S��\y��