�K%O�0���'nu-�O岵�ؘ�^F�eO�h"�]�����)R��1��6b�ذ$�7y��j�m������N��h?q���ys�{��)t�q�$���"Y�c�V�qЁ�F�́\�U��db�	�2#�Wq�����,�jl�C (1�]`
h�q���n��Kw�j�`�<ӫ�M�,C�A�(}N����u��ѧު8������ܢ�/HYX$��dU[i[/� �Z������l?SU�)�&Z��+Ab�^�H]�H����@���VqJ^kH �7
	�Pb$��X,�nDF���dZ�*Y ދ��f��m�9�Q��#h��T�VV�I�e���Fl���/2e�:��	����šg�t�16]Z��v-a9��-����1�P�6Y���ڸ��K�St�*���/�s��L�{KJK�K?�SE��O����5vaRɺp�ã�!�	�+���0�����٧i���� �\̦�6�X���x�v�sC��I�u�l��'"z�$�&b6P��.��Z+~��1S6����4�5	�L�E�PS�� ��P�����������K��m�	U�v����&ͦ�x{*㖣��^���ni,WU��CP�l�!�(�p��'��E
��R�i��A���kn&2�T@���85*������\ /�QI�2�c�b�|���LQ �3Ѵ�ױ<�X�{6[[��y���FԷǫ�K���?�N��F��   � ��u�&�k��Τ�d�&@���Y~J5����Ux- �58�6��۞�J'�#̥ȐT3�r0\�*'Ze+̞�T`�ӱ�׳�`�%�����5���,X�b�@���~��:��Z&�a��*�F��a�P|�n�u�c�:���ܦ� }�M*{k�1pVinԽ���(�9�;n��p;�7}c.띣�p:�����$�3wC��2?�n�"���M�J��g�zFd%�a���+8`��Bmމ�k�5�T[�h4� *%�`�k3	�Ҭf[�o��u���&�
���g�%�ĄԆ� ���H��1Mo�@�:{6q���:[G
(7�H�}�p��с#JQ��t�� U�j�l_�I�*٤����A�uq�4�0e�:"�mj�[)�����ͱ{���	���Ue����]V\�X�^�I�4���_�bQ��~�U���~G5k'� 4�|�ч|k��3Uř:�k҅�ɥn�:�%���E������|,�.����P+	5`?�C3҃<\���7q����2B��mea���E6d�7g�U�=f��垳E�si�!�s�	�RH$q}���Dإ?�H��S؉��P� ��q4�D���+��7�U/ae�Q\,��̲�l�<DG�d	L�$u�L�pH&�/x�
�bi:^�������R�1���R&���Q���p�/Dǜ��i��r�*ԉ��x����:[Jn��kr��
��!@!�d�yc� �f��{J����O�\1��L�̺>6}D�+��<"ͪ^<��V��ɪ�5ڊ]2�+Y�؄;:�C��30�l��3II��	]��'*-�loL���B��

֥U+�"tuiaRIv�Tc�|�2;��Yu<NEvj�F^�LT �Sէ�I����J�l߾��jc����]Jl���U۔Q�LϛtJ�v��YP��$�N�ݡ�͊ʑT�/8R���Fb���F/�~&��U�՗|���&���n��f��Ay��]�ɛ	��<�* ��*ͣCY�T{eu��`���]�+���zJ�o|�Š�$2n��)��m�DӦV���*oT��4�{|6Z$����)���R���i���Bv�ɱ�����; �z�qH��W
�\%�j99�6��fY@�sTK�K�i����T��u��^��'�]����ΜS�%�[�n+���-b�x�l8GG��`J}����`���=��2Z����:��R���,���?��%���������$L�%m��}z������9MO�c#�em�*��R>-��⛶����1�(y�8KYkh�K�">]��D:y�����Q�P����~�ڳ�0���LK_� b%�����>N%���ֈ`����T�&�ҢЦ�0��{4�I/��E��{��`�k�^:3:ZhN�����0*f�+8�^K[��|��@�H�>3�M7<a������N}��]�ʷ0 <>뀏�ѝ��MJ%*�6�h�A���a��g�D`4Ż�4
�Yx�m�aF�xA{����OǆVNP�F���6D@K���
n�
���ӂ�;�3�+@߯�����Xs^Y��ė-!E��������P��NxaE?Vc ����t�#��W�J	��n7��OA�'2�Q������1�YaD�a�nB�N�}0�y5�%�p��#�F��BE�;=��X��̩ץ�yb��O�6De/f�=6���h���� 8Ts�Y�v�����R��_�	j��v�k��;e�+s�N�P�0�:hP�D��   z ��-����3u�YR9�EB��B�b�B�[D<Pt�6�QL�T���:R�|${��!&"K�~�r������ꦓ���k�󎽵��{��3e���.�ުY�Kd��
lZ�|���$��`��t.�G$I�ӫ�z 4L'0˺��*�¾�Y?�|S���B���n�A��wF�YR���\���5����F��-L�/&RMxT��\�_xqY���D�<�N!�h�<aT��.���X���Z� �g���ei�T��ZάO���L�ˠ�\�2 �P��H�($HIHM�p w�`��jʮBNQ^��Om�o�V�F��m�v���e*@a���TH>�Bb-�_Zg.�%�.� �Yؐ���-�� r��m5yy:��0����=+󟮮U=ir�4��^˝���Z�pɏ�(���G�G.{�o� �[yM-)����6x-��/�n�������iIt-�[��I�-v��A]��2Z���z&�uA����J2�5�g6ZX$9�����iks��KC#F��B�Z����k*TP��^�;�-W�~��[��u:/�/��J+3`Y̤����|KB�-lK�7h�ۀ0�-#����`����g?$`h-&��#x�C��o1��\^�����n��5Dژ:C�ٯ���%��f�=x�(�{��l�c.66�5P�B�p3���{1�mU���=*V�s�4Y�ٻ�08^5z=����<�����2
x�����vl��9i�咶�k���V��w�!�%��ѿ)���q̔A+������F�ˉoT���htk^�&�8�Շ.wY1
�
�O�@�b�s#�����k-1�G[�i�����/��kI��H8�b�Y-�(N������������X֧ɕ�8�u�����YƆO���{�z�8,B/��D�
�YU,WN �8i���Hv'yB�f�C�9~���FW��^l�&�|��_G��]��^a��%xX�5�+��ɵ����%- !PRxV���.-��O� �׉p*������c���xΚ�ú����W�W>��_�^��ש0�P��Un�tBB�W��4�����&����Z�������#6 ��g��N�k�[�&ߤ���d}��   $u��U��D:0^7���!'䈝���.�֮6f0_�cf o���
�|I���#I�Cu��Ai�̞�e.�Yt�5��v�&(2���#^�W?	���S�y�bӈ�y3s�y(1vg�R�����W@������-'���_�apI���Ke��B|�ۍ��.���bj�D@��� K��� 9��{�b�R����� R�s�1�r��ik�ڿk��s�bl��r�K��70(�d�TIV	q���z�.��bj�C2����?� '���s��qlP5SA8Mx�0iU'A^VTy��-w� �z)w �iaW�JK�xc҄�+׹V�e���o\l��+p��6�I����_RREu�i�=������&�����ET�!�$-�ŧD�k�k�X�NH����6	�t�p�)7�AԌ))�3Ҥ�gC��f���F�}�'�b�jIK��)�����OS.'J�wň���V�]PBvt}/n��V,B$�V��������d�;dIx1��K�����2��_�|���8�٤���oc��ܤ��I�n�&�}�imr�kCp�˓�~���p�4	�b�0�%��5")�tm�K~��\<�N:������L�k;a'�F�KVc���5WR�Z� JcZ�l"9f����f{�!���heGK����:��*Y���
K�\���<߈i�Ĕ�߫��Mi'�g���K�/�im������j?D) <��J�y��D8z/����N��5�˼�w�h����U~�������'��z3q����\-�Y+�ȝߘ.0X��U�X��eHL���6�9�Ԕ���Ȋ+�F�qSSn�O�-��+��fX����%������o8�P)d�EЕsSؿ
��F%#!S[r�7��|.�+e����[�8DD��`����}v��vGn�⧈�V�^�|� �Q0��Ɓ4�+S>m�ai�P'51��X��5xO���]�?�Q�[L��_U�`��YSI�_x���5�z�q��.$괈OM'���g�ڈB��9�oT�Ww|;�l�<�;��g�+!ź=Ȧ�I����5���5�L/:�)'�A�6�T�U5VU����
��I�t�+y����ژ?���s$sxԋ�d�Er�:�âmu����k�����cr8�%%��D�)�����P�^�A5�yuo�Z����i���*���\��2�b�f�4�p�a����J���	&m�H�V,�0O{�����Sy��}4�R`���Yˀ%��g�2;���t���aU?�I���!x)���^��pU��e�7�\�O-�~[L�p�0B>͠&�jw�8#�/'�
�ĿG�b;K9:S�M���Iº����g+�	V%�~"�V���(�W�� �d��"?U˶��>�c�O0� 7X���������C����oL�P7�w�ƍ�+@�������F����_��t~�9�y*: ��i4�TYD4��՗L��u��z�F|W�Yą�=��<X2�jr�Udr�x�V���ß���*B�JSziZ\��sƹ�N��6�\�G<0<p`��%����r�<�/hx2ߦab�y��l(��|�	�Ĥm˃K)˰R�ta�߰�*��XE�|,������T(���Ş��<�j���Vk�o�~+�A]V؀B����I�Ռ^s`6�q��/��k<�%���%�3��R�'svjրV,�!�̵����������С�w�r^��u�3�	�?��*����D��q�:9j��y7=���$l/n�K�07��vCۻ�«���А^�>��LK�`��bѹ��3ӔV0ʟvI[�����t���	���Kx�e�p�i�2M<)eg�W)������+$� ��o��V�N5�/9��)�I_��{�5%2ԧ�ͅet�����V0�H�`l��01���{x��������g�O�Q�9���R�3!8I8S,g�� ,��&�:�i�f�t�b�����
v��	�09�ˇ�)]�@�~��R��3�N�ƓUr(t�)�*g�� ��*(m�e��߉1YQgUw� �!��sY�S�z�b���������ٵ��=����[k���y�l���(Z�g�f��L�� %�\��K���qg ,w4Q�B�G�|�!�N	8dB1�ϲ���5߁�jl���C�zS���Q�s�F5�X?���J��
����M�b��O��\-fc��22��ڪm�A�%~��\WA��������������l���xoIW'�J�����j��9�3�L:�v�+�bA��ʧ�޴�0K1�� |VOIF{/+�!nں[ʆ�op�V�ᵭ�]i���O5���tl��ٳYe�~�� ���N�k�
����o�10v��B��/�1��;ӣ2�j ��]�f�577
�KS�h�_��H~z��*tK4Ā�M�t�ϟ�j�q4T�m����ک�^2X,����з��Q��NT���w/vV	>6�S_p�g`��X�Ѐr����>�0^E|"�g�hR{��j���)�������ޡ�h��*�pbV��|�p$eM��[�t=x�ti+���������W��uXAT��p
����c�〼�^?�H-Q��ն�^4��I@	>E#nv0���&7��9(y�&�K}���&caR���U�>���RBo#g�z����y
	Ύ@S�)'s�u%	zv��c�5�Ia���RD�
�^,9tI>�-��4�f�#�=w����4� F	�ৄ	#��P<�\�s�+�Sfe>��Oj�搦�ݠ� ;B��Bh������6~�8�'K+B^,�7���v���s�d�|�a���
�]��xq�pX=��Щ@tJGte�����^p@�7{�Z���R��LiHu���;�v��uіؠ$��A<U��#����d��fiO�`̆�Z�S׮�G�� "A)�tD쨊/t/8��&��9�����ѲD��:���g�N�g|U?DL_��+�_�V�Mlz+�Q(}�*U��˶�S5�\�oH�H"b��	��f�T�Z�Rȸ��w��M7`���qeyiB��łH]/�Cz}zb� ��2��P��KZ*�_
�P�7sm4p�gA����� ��'+�CI-u+1|Ak����)W�/�\�b}6��;=N)�<�2UD-*'���8�;�����B%����3ݟp6.QE/��:�@�E�`3VB�-�#<�K"Z��c���~"`�r#sb�3��,,B�G�������o%y&j�*F ;ڣmt  zG�\=mAit�iO#�̪��&˸�B����OA�_z] 7%�������l���ʓҶ�B�+��xiTx��C34���H>|F��K��uT-��銀��''G�[�wA#k�`�o���lB]7naʠE7���{(�p�����Y�4U_�pv���T�(�r d[7��.u�/
���Did��U��T���4ٹ�T����!n؁�V�Z�ޡJ/�$�e�I6J�����==��Q�ĕ�`����~h�Y9�/x�L�9%�������U0"��I����w�0tBw��Х�
���o��p���)��2ę�B��rm�ю[�,c����k,U�a�u�=��
����m�޾�`�{+Jj����.��N	hpm�"W}���I	!�DӴNm3J{��+3�T�t�K�+�6N����'��eD� �Y����d�X��^��v݉X_#��;���u��^J:ƘW�"�Y�~��g�6�p���:0
D/�y��4��荿$��0&�/iS�~�(�WV0"��qg�8�l"�5r׾����g�.^U�z�|�=��_8u����o�ט>�l��D��l,�ӏ�k��G�%��bj=K5^W�(DM� um�1M�����v�1TY ������>����x#��hv�5ؙ��J��9�6����P�H;�lDO�pf<����fe�A��iZ�ڷ�Nb�BZg,بpLnoM�7��V�e��ٔr�����5�-�Q���ӟ���V�[爕����j��^cd�4iL`:@�˾��	^[F�`���Ѩ� ~��
�y��߼y�dP�d�O�1v�Q��H0���X#,P�0����vA�g.��4��m��󂸖"��
� X���j���e���#�`Bli޾��6������g{N���__�FG;�F��;^W-	���u&��/�I����:�͈��g�QH�G��O�̗�z���]�xNk.������E%pl�g�I��� �B@�L���3�ޔ�8V
T�$��׭L�������Q��b�ekڰ�#��Y���X?��-���9�"��V��M�ْ4�h�܁W�-��_�������{���UL&}���k����z��HR��.a���9泺���V�5������ė��O�e o���ǎ�