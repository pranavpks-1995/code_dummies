�qy�p��Lx.�V�Q8�\��u�ޑ��i��ϗ��u��͛�v�oϻv���e�,O>V�˖�����ӀW�v8gy9��6��{ׯ��6�b���%&M��5ZE#��a���������`I ��e�3]Rތ��a@��čy���բ�dį�t���KU�=���	�}�2��ԨنR�ڃ��x���"�#ͱˇ��Ø]�(	:�'�Lx6��]�YQ&~��i�2'?~Z9�k�����.4��~i�K�<�T��	�>Υ��ȢC������ן�+T	a�Y��'I���׏�K t~�.��X� B��k��c����pY6w]n��}���d��J��K5��7����*Ed���q���0��W��Q�]-���b궵6criL{�G�3~� �.R��IR�����m[�~S!1�D��	w������2"�dz �ΛY��c��
�NBvSAs��v0X�8N��a�ph���i oT#��\�n�H*wCNmg�����:��`}tu0"� ����Bi�^B��G`Jh��� ڳQ־�i��?�~
�T7�oZ�	Ye��8�Z%��Ph�>g���՛�4d&ύ┬�������Nt�1�~u�Ϯ�?�!��������	����UQ����P<�;|%Zu�`���t�2	3@=t����M��+j�[m�W�͟	����v��I��@iy����e�/`p�������Q\$��+�#Wy�Z�H+/�Ń�ӌI)��i�M�g��{�'�{&w�Ӷq�FVӂs�31l�7�}�T2���Kއ�@*̢�.�	�z*�cO�|K5�q�Ɨg���(���MAy�o��ʒ^![�31���\A��}�x&�%P�(:䙝ŹefR�;�U��q� "���*A��:E"�=pQ�3��v�%�c��Qd�&�,�J�%�T&���O.6$W�F��8�L/�_}�&��1",|�J�ڟrT���H�yO� ����Ӏ���=�xN"�wG��\8��O�r��v2DP������@,j	�|kԧ��]�kz�>'������^��F�3 ���mŅ�f9�S
�O���!4-`z:�w��;F�q���5l��t<���������6�������y�4M��Y�K��B�(s���5��UZ
����< ��C��S�_J�U���ىP����#�p#t˷�n��N˖;x�U�}������Q��G�.�!�M�]Lj]�ֹ���!�enn1ķ6~_�ȴI��6��"��È�/^�k`��(�8+�g�n����������5Ώ1��>��P�X`�|�"�G�����Ju�˦a��n;�+�E�y�)#��<�/����{�������-,bǧb���'�����a3*�6��B\�w�&�aݯk�ˏ=�3������)̇�@��G��wb�J�5@jFE��n|L�U{ӕk&�ϱ��%�iɹ�cT�B��b��i��h�⇅����Qo"4g�Pl��F�Q%�`2�R��z��u+�8����3��[��5�D��1�� �FB�Á�DZ��|���3�H�r���挍P�p讇{�y�4*J�X��U�y�靂��.aIx���טO��)�r>t��W���~lh����4*�)[.�~B�vl뙈(h��)I��<�w*��A��&V��1��gEq�W9�5��(XY�sv=�ٿ���L�%�i#~^r�ܽ���]��������)�����?�l����J<p{Bi8xa�^��g��I>�N�|N�R;0�N4ay��{�QnM��c�y;��z�7r�լ
g�D�z=&��(վkR� 8V)v�@l"�м�PA���v%-�F��m�D�QHZ8�#;�EX|�x��X�ܖ��E�M�m'^��g�ȟ	�'�:$���&�t���k�=�ӊ������m��ބKK5���ۀ��*.v�솂�i�<���K�ߞ�<�Wа��;�����1�t��ḡ�����5N]�/{G�~u����<�����j%BM�tM�0�x�̦@�����`"��	��$���u4�o�a��]�
O�4!���c����K����֖;�;p\�����c���N�T3������u$'��g'Ђ�\���}+�QN�����y~���H�o�7d����������#N_aS[%�u!���q��R�|�K^2t�k���R@�[�8�Di_���s�c���ee��&��\)�
�>�u�#��DCp�ҤE��BZ�@���^�R��;r����a䇂H�	}cV�E"'XAq��:e '�
��]�it��V[���Hߗ����IA����Bv�������H���X�(��&�:��`΃��5�~+��:2�["Kd�-�nO�t��\ NK��%���"1�5�̦�gk�����27�J�A�8�Bo��무�r�cW@y���H����:���n4g�ޘR��&�f�SJ�'%�k��E��Xm���#�z��
�
qZH��h��8@�{d�?!����P�f��j�g�ZOwW��n�Z��z�Jm�^�:"��C���Xze$m8ù
jC?���I�>���&��#��.�ܲIܣ���sx �f�єD78x�_|mU��ڸa�"��uk�����g�%�|��?��z��t�6&4򿷦B醏=�P����ǖVk�[F�f@���H���GI~��73��%p$��0@��S�շ�����E��-�2�4����c��F����x�W4�v�m$tE���Y�vm
���-��z�K}��ڼ��7��%d�7�۴nך_#���'S�;�9q+�8���a=q�UéN.N"�����"Q�oj�P�����P�kh|xC��}����Ǩ_���KS"��y��e뫊1�KX��2]1a򺥶D�ɔ�������ۿݛ�@p��c�H�����@C9ĵ��?���"߸���(JV(r����x�P%��:f��P4��k
�������� r!7yoѠ\�z���&e�W�VY%����-Fֱ����#�?�+��i���m�X�#s����=�{����6IK\���!C�u��k��p���;]R�?8<T#*��	��|<6K7��yz�9fS7��0=� r�g���\�"wB�7� �\���Y'�/��L[�4hZ9ш^���'%b�2mɦZ<4�7��wu =m9��<ui�zB�f(������HJcy�y�M��&��hO�<5�<K|0�LB�2�I��~�o�x���D3Y��|P�Х�!'��~�v��J%�_��e#�B��ne s4�3�T:���F�0L��xޭC%ӈGOO�O�c�ٞ�:���b����j����eE �3��4�H����c:nV˩�Ou�>��ӧ��ü�	�xQظ�1�����|V�ֈ`FzSl���⤫��Fl<Э㞆t!�ir�t0^��W'��g;ێ��#���0Y	n��/��ݼ�/�R���b(���������ݽ5Lo}z�h��!���.�K^� �HQ(9�X�|��g��U�f���l�;��m��RdU��8�����yv.˻gY�Z��\E�A�*�������l�OU�pV��v��K��&���Q�Ӯ|��g�����L\M�F�L�s:��$&����ߣ�0���E���:�3#��퉺)$�?�eE2P���E�J��1삟���B� ��q'�U+Z�8�J�&Yy��[�?�5>ԏ��r����婬·�ީ�ֽ;P�;�S\-@����P�y�m���X���D��@��-���0JL6�?'�}����f�^E��W)��6�-��W⟽+Xz~���.Q�W�)e<��-��۫��L�7�k�A��*���\W�Γ�!����:�hDJɀ!��BU�<V���P�XW�arɹ����e<��z`���;~2�>�������(�$��	Df�Ow�Pk<���Y��l�o
pb������Cde�Z(ʄH�x���F��#��>��η�c`�X�PIQ���r�$5>��lQ��R�KQ�ɻ��6�|󖟭�����N	�J��c`<��s�;�k��}����+S�ɠ	c��4mG���Ax{���ԍ	���5�Q,�h9��=R�A�%����JGLG���UI��+<�*�O�][+�%(Q��fD�F	�N��x"�j�N� �������{�����yʯ�_��ɵ�B�#07��2�)�N\�[����/sm/�y���3�+,����7�x�N��r��}H΍E|�ڈ�=�{z�a8�������E��\7�B�GJ���C�?W�� ��h~��xt�H����2[{��R�y-�ó���w�M�ɍp��v8]�A��"�=g;�iRZ:�W�����
�z��W� ��G"%��G���.���	�����ʐ1���}��Kw��ĝ��l#�\�sS���AN��|�V�����޶ˀK�踈���sA�km���+ҵ/��ϊE��N�S���z�heV�h��nn����ZӇ���ѪRVZ+�[CXz:	�"��ٝk�վ����������G<��Ac=������0�-wfF�e�]�0D?m�������ݥ��RY ](��$��F'0y���d��;�����/����n���=��]��΄�Ӏ���{�1 1a�3�O��s�V]�%q2 *�F��P��;��a����>��6��!��5��^��Zi �Y���T�{o?	��J��-��?H�׉�%�^����L�yZ�2�<�ѩL��R��6��H��'�:��b�90N��6��L���lC&��s1�N^���mJ`'i`��Լ{�%g��ܸ���.;P���A�K�R~�j��<������0P78�f���P�Y|
E���Ş�$dL(C��ؼ[��t�,���~�ܷ����.�`_cI� ����j=ܯ��-��/*���q��ׂe1�r��bQjX�Q��[��7��qڷd�;�S��漩``�?���	��G�w�F@}r!���7���>є؂�diW=6м0PW9ő��tT�`����NH��E�#
�v�6~1���a�F;vD���61�0��r>��f�$��i��'�;S�@ң.���f��O�h��6�p{}�����������⮵Lm͑���I�C�*q�i�+�W���1��3D��~��}��l�	�f1��Z��4L
o�lD���-9=T1�>˝_�E�zb�	��]�ǵ,�����_=b|��m��]*�F��g���k��yVIN$-g�d>˹��}����gX��	��[����!|v���1��3�Lct�z��{i^�ٶ�5[�к���-@�>��X�g�q�"������TUoac���)b*�	Pe��X$D,#�HC��\���&��7��@(�����(ʊ-,h�7�#C)n���p�!��`l�a��d��։�D�9!70��0״,��2�Qմkt�7y=����OW��ʣ�qc�D#hm�|���D�ϫ�Bh���6��@�D+ ��LX��5�*kO�ց�hԲ�8��~��&��-��p[����a)yĸ��2W�W
��Bs����-@��)�jcc�d����8͏��)�&�|���J���A�*�v�s-��E(�lw�WQm����[���7���1wq{ӝrA��j�#���n��eFy�%���1S>��xMH5�42�)�
�:x/Q��W�](ZJ�H�~�Ǥ�h���y�w�?��]^x��@
��Rdm�����t�zC��dZ�(���x͏hΤ��)�{c�%ۡ2v�e����M�rZ�,���Bh?�J��V�_A�E����P�z/E�|#)ߥ��#v;X
d׼��.?�z�?H��K+�3�y�ae�)�y�J���اԪ3J5\�&'m�tk�ײ��MK|��x�7����� ����Ts��a�˗��� �8
u)��/�K	R�ve�>l��#��߻��5�(KP߹l��@j��������&�?3�+N�
uk���� �a�=g��\�A�.R�gjz  ~=BiV�o�Y�bQ�k�g�^��p�i("HUA�����W N�f�Իq8�!�EIݤy��Ҋ$�φٗ�<�&�j�(N!�(J���C�,#5Q=��}.�k�:�{�ZU>8�>����Z|�;���\�w y볪%/1�Hvix3qr�����ݕ< {ݎ|��d���ٟr��s��hR� �:�z��>���W1�TԍRѴS:���)Kv4��R���ѳ�qE2��#���x�q��V�X)���s
̲.�C؜�9&,�ẃg�$�ע�C0��R]a ��]Yw�_S{"�菾�~��`�j
���VH��~q�A�L|�4-B!}	}�~��+����$$��gIZ2���%���[�i}�y�_�ܯ��)�E��O�K:M���(��W=�H<��D�)���t��<:��B]'�O<;��e[{�u�M�vO😵�j/�Q�
N;��,0?��/���rԷ�@'6>��|���)A����d�طh�%u�i�{�u�<�Sh�R��:�@�Y��^B�'�Ӱ�
���2�BdWb���+Q[z�{Ө9r��\O��`�~K㽳�M�������Bn�B2��L��$lȢ~9̹���)�-,�<��|4j�j�Z0���$��#�Rh��
X�η4է���8�2Rû�o:g�����f���y^�VY��+�ȃ����<s�a� ���y1��R=�kɚ=���9� �嚸��P^/��2�t�Wz�z�JOM����0#�b�����W65Z`H��w�Jc�X8<���f=���FU2a�x0���E�p��2������t��a�t���1�M8���ۡ<������d����4)~�ﶦ3X6S}~�ٻ�=����4����"s 4E�]"k��q.��a+\���8྿=*��q/	�4��� Mb4�����n���k��%J�1n_�������&F�V�W����|��۫�*!���x���i��Ӓ�:�~��R�V
q]&�r/Rq娿 ��>Ѽx�����1?$�Zb?^�5����->���Z�P�����ت���`���p�J�g��, Kx 9x��}V�\ԯ��e�}���}В	� L��b]�9[�8�~^�^��cP�ށ�c$�3�,�FF-�
�rA s��!P$V>\�����n>8�lۣY�~e�S�s	�2����&|&�q�Kl%*2����z'��a�MF.��I���5ټ`��-h8T�E�Hg���{�!�ߧ��vu��	[|��Y���y��3IhB�cz�Um������Q�(-����堄��L ��B�����9��m	­�5݁�xs���/���H�ug�T�2������eߨc��\��q���~G�PO3�9Nr5�["�*fgkx1' �X@U� ��8]�e ���_����,l�H���L;�, g��`e�Mu���T1��+V�b���	�.�j��^������=���?σT{�`!R��u�B]��8)��V�0W���Rs���d�	ܰD�������F�pYC��0]���H��tk$p�&i�*��I�J{e��$ߟƏ��e�A�Lu��1��A�"r��֎&$fo���UM;vn�a���KkϸC���<�0�*�����y��7� �#DƟ��g�u�7�
�u�8��;@+o6I��妾2�=����J�|�U�ނ���G�F'Q��b��n����F��-6tm���2q�D*j-Jl����	oՙ&�4n�+�.�Xx��(���ρ+U���T�M4�\a}�T2_���'"�i-[Ր��1�4]�gx�Ś�G�7�W����-[g��>m��W��
���s�(���p�)f�W�)(К8��<��;���R�S8Ϭ���:�7�Z|�4���U5��hCA�����c�B�q�@�Cv��Q'�Br�D|�=Ua��%�9rl��Do���T�Pl;�?�3�%�,f�5����bK!~��4�"/�]7H/cc���a��9�Fvy�w+�D 	>1�WX�L��o_�=�D�NS��"���Z����Ej��U,�c�Tav�c3$���+`ɓ�2
�}@F���f7 ���\$�	m���������?-���g$0��E]_í{Q2�(��,������ �I��!x����vH�iL��>�5J�U�#���h��U쮔�o1�:'�����1HCE{rL=��+�I���u�������gWZ�Ư�<�2T�4�`N��*�lט�6;F)��yI�kj��� @MZ��'�5eH�H�<a�P�����/��A��6��#a0�Qk�U>���K$0u��zZ���=�+�iݼD�"5L�K�_���;�%�w����-e�CB�!M_��yr�|����-�pƛgej쿙>u�+!<f��2��g���sG{����Бu`��YA�EfRz
��Vr�H�Fй����~�^�����w�9��C�8�)&t�����	�uǜ��z���eD�)���dK���M�Ǎ�t�"�ePFo�)(�FŴ�D>�H��_�(-�
ed��C|0~2Cj����.ׇ���.���0Q�D��,r�>�j4Z9�N��Q<	�b�l�ǩm�%������'J���vh���*-K���N�V�_��*�)��fx�U��{'���nq*\:j
��rY*B�2	�>��<�$�0�0���=b4gΆ��Z��$��/G��$�U��k*���_��kmE���=�\�2�y���)��]�A��Z��^w��E ~.����iD��GK�6�INs^	/��Q�9b^h7^��U�Tw�8ݓ�?�
R$��ȲN"=N9����$c)����9	Y��H��lЙ����zZ�_�7����5�� �,��JlEB�?�
5!^񝼱C�� q�~an�++ݯ�L��VA��j�ڪX���(ʆa$�fNf�'�38�>�v��^��VT��}��3�.uJ�m��0"��n��z���_0�Q�{Zd~{����r�I��>�ȝ,aӣ��$�}O�si�6�V���"�⌹l��[FWr��/�
�nf�w����KSY���ܐ�`r?pOOB� |������|CY��4=����Ǣ�XW��l��[���y8ϙ�U������4 '��7���OyyfUd����Jq��B����K%����Ҟ�Ȟ�
�]թ��oe�3�L�8��F�7U����ns�f-������ X�	Ｂ��'�D�,n@��z_O%N�jTj�E��bmjy9{[\8�0�3�ʂ��J�:���t�Co;g�%�dM"S��_����_ނP97l���z��"����i��1���׋���G �ů���Q2<�W�aJ rj�ۘB��u�f���vlQ�T��=�'��z��(B���QgTM*BU����Jc��!G�,��t#a�4���0,��k��ѐ�;nhA/l�L���>��/5�U��%=��ݲ�!�r|�;,C�4��O4��3�h��W$�P'�y��l�>�@��$�s�&�M��I�wP����'�L����Fn5>�ަ]��Ei���)������s�=70Jc|�1�3\���ǝ�������	���GGI�G �FN�BlU���I�,z�kAa�j�KY�o�����Ē�-B�np��ѓ�U����adX�*����5��������|�]U�x��W����>�\w�&tT���l\��)6�'��
�h�&�٩ # Ek���{v����c*跟*�C[�{��7�q�:���k����ח��� h\���p�1�]����zzW�r������Ąs�%�.�x����s������]W�����~��>����s3@�m��8�`ۧ���֏�y�5�I�	fP��kfewԹ��h#ܩ�L��Y�	���kbsE�w�ut}c�a0�ޕ�j+`_A�I%}�\�HT>c]ދ+N������2z��OX�y{d��2�������1��ƃ;��1	��ŋZ�������ŷ�������z7>��QvB�R�Ӹ�|�i������V�mL7�j��t)�=�&3�;-�*~�,�Z;�M�f��cu:��j�i�a3�~��@�B0$�VV��h��g7Ȋ����1�Ԟu��うX���g$`�G[��Q�}����c�S}����7�Q�tlp��п��y�қ�lodc]�*Ԅ���瑼�瘢|���T�ǃ:�q����o���-�.��Lu�<�ؿ��n�� ���n�n����$�} 槌�jN"��*S������3��w��f�]�Pƒ?̌��Q�+^���T�7j�C��lƸ���i���������E�=����V <ϴ�=#��A�����j����;��a���ﻐ�)^�(
`砊�mĆC��i-ɗ�At�M�`l���Q~�?�7�L�	>��Y��aDґ�#�:1b��!
��_v�KS� sW7W��a�B��3�+,�����-�������^���n�f�z?���i��3�r.��qy��y�e4w}l�Hʯ�~�T�m�XɎgVδ�irYo8ϚZ�ϩ�� ��Jb_Y�G4+���AP�H&�R��~����'� +]�4��!`N/� c��͒�M���HN��� {jt���:��[�ʼ�����K���{M�sAo��}v0�B1<;N���3�+[а�?n���4�}�a�K�P�Grp �>m�O�x5*��Ő�o���x�@7r���A��W��Ǳ�8[7�M��@(1���1��X�8L�����ʡ>�eEL�^Ɍ�W�j�܁�r�ͺ��ZJ���QJ��Y:���<�0�[�s`��:���g�X��㽗p�@�-�Dk������&��#���Un�oJh�ֹ�����}�����!څv���)zs���?q��Ң��	 ��ǭ�vm��X*h�plR����{��,�Q�,����T��c�F�eh}�dݼ������]�7Mss�5���('?�Z�JN��D�%���S���ś7�>`|���!ҫx�%g!��.4L�9��oH�K����_?�Ac ���behrO��񆈄:N�\}��o4�+��k����j�����9z�i����0`j*& �6`b�i�ڠ���`���g��W�� ��'���U|{�y�/\��S��ޖ�
_^�k"mEO�]#�������oL�[y�V�Е��� @��Y���jT��ے�n�s��r�����d�6I�4�0�j���64��5N�) t�?
r:C9��m�)���){`�g��]����&9�d�o�	���(㦵#�l�ɓ��^�@V f�?��"3{x��;��15g�	!���䁙ڪEn��w�L��\��J���u��^pU9�6s �ҳm����vbi8�Ƅ��c{���"�y\V��������5�O�3.D>���"���?-����+Qg2��*j�XM}����\ (�-;tP�θ&K��?�ZCE���� ��}#�3TF�W�8к֬�t�<%���]�f`��"2�=׳�6؆�}H�����;F�^���������&��E^m?��Y2�vgM"�_�.��y��]�w,F�����Èz�XLS�}\@Q�! ��+��P�h�(D�S�	)�ٖ�
j0h����$��B�ԗ�M_�x�
�O�Zrs���*�n8�N&3�U�W�EIC��`��*p�Cu��_8��&Ǉ�<G�8��w��>Y��æ�Bu�^>.^��)����:���q��))9�D������v(~+�77��nu��9��k��;���*�3�%��fF�2tD� [�������� ����%`��ZH�[ѕ�׳�!��G�/xf��~�K~U�k��]j�a!~l�z�%��V7�%�UO�LE�IZ:���1��H���K����@lx6��O��e��<e�|%���K#T!_�e��a�d>2�:Z���i: �H��Ĩ�B��4�*�?���d��
'���G@�)I��v(@
�p�҂�Q<�:�`KPf��J����Y8��W���0d�*5e�+4 Y���!��<o&8�d�u2׋`$F#2�,1Sw`��'�9���q����>c2��o�R7���uQ6��gt�x�ǺF��3Y��QD��KC��ݓ 2�|�r���$?p@��T����8(��*����,tV��5=����;��2N�	D�����S�Z���>�a�w%��6�N�Gב:"{�G'�D�r��ťSm/���>�L[�n���sǯ=�WW��a���"���T�D\�ߨ�<��,�����5IԷ�F�I�I|�@R�Q����z����EJ^_���9��g�Q庒KL*����������zo���p����]VA�vmد�mm�Uj0����7w�4��A0�L�~6�E7f�?���g��e��շ����M��_�lX{�	΢��Sj~��`��$�^�����Wt5�j>'HUWً���*�ݼ?�P7Q��[�eR��>���5�-Q��C�pC�9�ǩLC~'�%T�U�F\9���N��}39����m?
��d�e3�đ�B�%�0*`�[��EƘ�vBx�q�<*�gU!���	�[e `0�! ��`��[� �_��hAZ���C$;���}�bA=D�|��t,+K��y)�J՜�	��$�P�/T��WGȹ��r������z+�8�'K�p�9E�I�Y/=�8a�yI��T؀�����>����%�e��h�6<�u$S���ٕ�{�j*���r��5'A����gW4�{Ys�`�'g}{r�t��~�ںL��@}>q�P��7�Ї%3��V*^�/!4-�&}گ��ڧ&m$9s���2�γ_2C���Y��+���7k�eF���l {�Q!���m�Վ��Z/k��[k#o���o�	�X��S�\ϥ�A ����p�"p�B\/&�/��6����2|*1����{
��^�[�L�%���{�"��7�vHpw���1�FCN~٥hA�>��JT�)N�n#"���k� y �;�O7����#+������=���\y6�����)�����:�n>��*��TB�[�73�2$H��Y~M�΀J��#DV�H��Z�y��l(/�̶f�l��#�ǂGu�� i�"�
4�z�5��4x>�JMy������rW ����p`-�_ ��pϋ$W�k/1��%^i��e����o�H�ǵ�@�\�i���,�jW_�=��x$qѷ͍�$~JD6�.��@=�����+�{W���X̟^�{�_���,ծp�*em�N���ַI� X�a�G:�t�����Y�Ğ��;_�k�v��:Ok��OAޚ� e�0��A3#"���������o��U�v��i{��l	� ��ї�3���.�����������)o���2Q����q�?GA��t"�ЍAK�8��T��c�#�s�������NH��ҩ�>z;���S�p����%��=�2����T*}�k�w�\��V"���n��4T]"��4��
h����5��$ʅ(��oZ!7���q��i����P�	Yw��l�T��HX M/EΓ�X��aҜ>a]�#��-Ƽ��9(�8�׭p���ى�yĎ�"ɘ�j��p'���Ǩ|�V���9|�o.�ɽ���X�%ю���UY���JC>�rl�[kƙ8�֚��}������ΩS�!��mC�ć�9Tn+��v]/a4>�o>�ݱ�c���g�9͒j�j�SzM���D'�f�G���y�e����ۙfE��*i�X|�O��!niW�Ԇm��� U��6[]��Di��}�sbo95�'�Dɍ���w39rZ��tw�T�^����X���
���] EJ���ຮ��H�T	t��xD��B9~\�eJY,m�j;�|�^�5�c�V�BX�M���8���@{�w���o&XSǎ�����!���^y����V�v���`iZ�#��x�	T������</M�~2�p�ڄ���c"S%+Q�> 69N�v�_&�4[,��ׅрe��aV��ۗ�����q���~��2���2�a�����r��S�zd�=tU5̍B��"�TD[�&*�E�اp��2&J��~����=v8���z#��:5��(�#f�{�F���`'4�էwtȫ��',z��<i>��V�q��^E||�焁({���������E��K�Bb�_%��k~g��� ����#��Pؐ,�!T��;brE�.�#gM�#����S�$�wIS��珣wE���W�3߳.��z��D���E����S�Ci��E�� ��������!�����U<e�n@un�V4������늈	]Ln��@e�"�KZsdD��
���n���E�����$L�bZ�B�/�R�#��� �g= ې��z�8�@��i'�)� �S�*��Ds�L���`��" �60�X}.��/ζ�� ^�U��YPPv����L��\E�� !��������fh���
�{f���k.�⡬V�S뿃t _:����|p���p��2��1;��D�B�|���׍����h�3!�D��r*� ���D�)�� �5`Z)Y�q�7�2�a��~JqvB�X$O㲮� ��XS�i� u0]B�P6�
��D�����p!��5.nr۳���֯�[�p ����i����`7�N�@��T�?��i2��B�M�����Q�& ���H	33�����V�9���\�UxԢ��C`	�A0R7��'`�� "�Ew~=eʗ�9?�(é,�����X�~7K1z�f
=N��3��c�)�I�M���!UQXU�G<,i��!��`�6s[` 6���.����I�A"[E7짾#����x��u ��;5�0��@-�<J�²��ji�����qSbZ�9�m~�.�����p���x.�
��V�� AB|�{�0񷑫��Nu4ƌ[8E��L�֌n"�������s����6�P^xje��u��!UR%��<�- !���#����ـi�.׬�q�R�аL���"^)-۬��T�aHY� l��W��H{?�AH�J��! N�($"Y#U�W�%V�b�+�#hP�`�.�,���ۚӥ�̝�|�=�o��2k���R�nv��4)����`��uޓ�����mwuUUR�%o�I*�{A !�M F ��P�(��M^��;�(�(���o�
Z���ZH����.+9����p�;!U���8L�D�r�ɺ@�i3
6�&T�P�;�O�jv���5 /�k'��3����r�npH�T��v}��eu�>�a`X�LX
� P7�hꪝ�wq���;�J��  p!��$/��0� q����t��<xʆ��Vk!�0�n��HꢔG)�s�y����F���Y�[ܑk��UpZa�#H^ē�| � (�g�E :�� c�'���gDY��o���uws+zڤU�8
w�?�"��<�, 4X�["!5��7��*�%f[[��k2 p!��Hf-���ߚ؋��2#��$t!�T��lb�"Ma�-���^X�c+,+�:'5ͳ��2y�J4O�Ђ
zWP��R����'�� ՝���9f��W�<�9kٍ��' Ż�mK�b��WYn yfRv��{��Uv����.着�Č�V��VꙊ ��Hs� �   kҩK�c��#���%!��F!x�	2�VF;�e\A�/)CCUW�O>i��<�R�;�Ʃ���g��1���x�a8X<��a��´��2J�}��b��(�6��yL;X����)f�/�C���Z����3g� q ��Mg���i�f��@�m+���Ѭ҇e�r���`&�jN
��P�U�Y�3^�������!vd&#>-k}�x��:|cV�u��)Ώ3��&��( j��Q;�אlJ�O���>�#HGy�M�ކ[���	��0�e���� '*��o)2�����Kb�����ZT�|M��br �WV���L��MiUi������g_u<�O�鍆o�ˉ��*N�&�����i>�5}��=_����(��[$�wG&#2�^	j`�&`�b�Cu^ȣ>r毖Y�6��zS)q`����v?ŖZ(
q�q��9)��>bwj~s��ؕ�4�5�t����<��=?���l���vt�W �@0��Lc��������6~�A�D�S��d�e���OW����J\5���G�/�ͫ<z0k�չ!�.S��&�>hD��@�fj�.@��r������劶 G@�H�����FC^T~�Zn���&0�>ڐ���x�)���4E���
��ʽè��5(��G��:��Υ��U��C�b.�sy��uԥh������ĥ�D����X�^,{>���l~:��K6�z+�x�_R������i���bc��;�E���N)u+�����{n\�_j���Z�B����Iむ����u�4 i��/�nV�od���qȶli��峱�e|#H�j����Ҫns^:�R���=��,��l�L���;A]yPX�E��]z��]�i��;�������c^���z6`Ul����ڊUWeN5����p��=�5��X/s>��=\:���k�፿� ��3��׾��
S��4�L�x����Q�Gњi�I�����]������r]Ͼ��%y6�#�P�n��h�l�fC�.w<ϿцwmJ��eG�1=D�gތ�\���kw,����baD�"P�@IvM.$-���=M}?�j�����=#�����;.]ʡMGj<�ܖ}�!�p����/�1�{�d��$e6_�}<�cBx���5
 �i��v�c
�o��%�ٲ���&f�#/�]���:�a�dV(��D�#a��!��C(�f��O�4�lr�t�X��=��l|I��.�1�� �A��v��`��D�#Q��+$�Bܕ�>%`��������]�2�U�f1�<�i
Q��Y��?���N�o�H���� `�����W��0JHn�3���c|��D����Rv>X�r^7��c��7��~%�8+F����;Tc�K���~�;��y��n�[e]�P�v��$�l]��{����^�����Yǜd)�M����7�
p ���Aj1�c�;&�~vǏ	"W$���j�=5���/M�#4?7�-���g��F� �t�Kޅ_�����8�$����H����ǤBȀ��(�.�`�[�b?M;-���}�Υs�2^��us͎{��:���_�T�R>���R9:	���-S�^�6�@��|#��/�ݨh$����������Kk�s8=f�f�ۭ�s�tx��e3/� ��/=ݶ��-�	�$*�q8��l<C0n�3j�����ĸ(W�����G����pR����k��4�G]@;Q�=7+0jj��9��rڬ�Oya�~Z�F�^aLZ|��ҙP�;۠��Vۮ�k�ڱ��k��Gt6��{5r'3�{*�\��oW�g���� ��� z��K�}<���k�W��bt
�W x!:Ѓ6��O!�Kر�Y��/�2��ݘ	�蒉��C~�CT�Rn���W���5����	���Ons[�E�ٗ�:F�����iA#<����+�GqpejQ�K�	�����7��-Q>���I�A����e��VY��µ��ؗF��]��K�(�/*
�ZZ���ͣ0����;�T`F2F���4�M�[R)���)��:�Epr)9���@�Th%�9��I��6���&�ќ�g����w��ʺ��ܮPP�!�������8���>�Pl5�e�G�JY	�9>ҳ� T��A�� }  ��d�xc��RF�#Dd@x�r&�_�	��ۑ{�&
�9g'����1J$�l(	��U*�خ-ŉ��B��>v���-m,0{����+���XRl߿�F��{p��u�