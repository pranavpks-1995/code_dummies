'T���Iޛ`��3$�z'Î@R����wq9 \b�eG���.̬���G1"���?2�F�]�UI��}l_c��;��$��,�A�/�@�	:�9���ZO���bp�1�5�/3�C�BҐN���~EiJ�=eH�/�ｭ��5�u�ٷKf�����ew��h��j�6M/�Q�M6��d�C�Z;T.K��V9eܤh�qa�Nۇ:�3�>����̋8�Ɍ\E͈�ey	`Τ�<�8"��͘w\H��Љ��<�bO�vgr��e��Bk��<R����jU�P/c��%�Ȏb��!�s��<�Cl/l�Ȁs�/N� ���� �I����� 	<����a~f�,	v�JYm��j(�M[��1׽�4f�!�gqIz��l��4��U���pf����eKW�հ��=Z���A�A9����F�v�����PKe����
������Ë��
��3�H\� Q}"�D�[�L� �b�vW�
���z��Y�Ǒ%����8[P��֑fA!U���������٣!�d";��/ёJ����Y�B��0T)-v_���圣Y����;�8�6�U6El�m	���Z_Ͼ���v�P�(Ҿ�9����C�ۤ��S)���+���,�����Q��;���Y~y�'~�����������V�����!�L��fܷ��B᳾Kظc��7գ��Ց�d��2..��Ԍy��UR����ob��O�1~��Bn|��8C�9�ƣ{Gz�w6т�����w߃^�a=҅N�j��_���	�Н�4͑�[o��P��M��q�(-w�c6qqF����2��[�h>Z{y£N�>ܤ�d�9z�j�R����*fؑi���΋F��V9D�2^�.1��IN }�����L$F�!ɩ)a�N���Su������Fg���A��R�p@NBY�q֠�0$��h��rt�ID����A�Wr�J�S��ٙ0Y߹�Ų�%��PY֏��п��zk�9��{�,�{�����vY-�śa�ek�;DE� ����4Q�8@V���rޠ�;�(e��$Ys����N=����e9����.!һɐ�F/�\��mG���Gu!��ۓ�>r,Y���m���ʭ}����z}Ê����$��r��O)��UI� ���=�/�ʀph�<lJ[qv;�E˴��3�u�e�}l�T�Ď���N�9'5�OZ�g��A,�
��Г�������c�4r_h�'O� ����:v�v�z�?��v�j�C�J�\���vG9��̘-���!��܉O9��?�e�f� �0(����E~Pԉ2��E5�:�%�S{�+v�J��)\��h���ɟ�iulʃ��pi�K^���'Y̜�_����ٷ.�;0���)��-�+�$żC08��^��(mt�ޫ kK������Xܖs5=t�3b:�ݕmp��r2	�jjs�L���l6��:�����5���TGV�������«���ŲdaC�р�?��8Q�D$�D��p�^��9�p�}@xb?x��"<&Y� i>1AC:G��,�{"F���7M�?���R
�u���tc7�(�UkD\���5'��]2�y��H���X���7>�§um�Hh�R/y9�&D��"�<��t��u�>@5�u�����ܹ�c�fmW5�P}�\�����b��Vp$�i�Fi?�c6��K�Ck܁��[K#�
�{h�^*���4%xX�
�^�u�9Qؐ�my�@7(�3CU�/6l^�E���r�Y��1�d�_��
�^]��(ð�C��&  ��"'R��c�N9(`2�@���zs���d=y��٭ [��Ἃ��;�4_(-^UH���-�W�m�,��U����G�(c&o&���;u6o<+���t�|��Ŗ*;zjj����v��V�qV�{aҚ%�J�_�_#�Yx�ܗ��x���DZ�^��,�Fd�e̠5��9t��H�4�@�:�_H��!��|l%�@�y�&���FC���ܛ�w�U�f�+�?�#�Q|w�RЏ��J��:��D�Jh��n�^{E�݌�g���ײч �����������"��	��f�1pP�5���
�1;5ē.��c��}�ߣ�J`��Ҩ���;р���3	yV�&������zCQ�v���,��������ן�6��xF��f/|��gY���'�y��'Kv�H�ʧ'�V�Ͽ]'X�.e@vvݦ�4�s	#��,�����3LDVlX�t�$��e�Qb�4'x��><p��j�#��t�|�̀�[H�әFɌM���1
��Bx�4�z��bb�r�K�lD\��k�:E:bh�Ik���n�|��g(�к�fOw��
4{U����,ׇr���,��\�i1�@Ǚ��r��b�J�������$���4!�}P���%�awvZ~���֚+�Luܻ42Nw�|,O��{!}�ج&{2��þ:r�6	��HM��}�W.3�����b��H���q,�psʧ�T���KH��ԩ#�SF��X�ɳ�WͺL"grz��Mc����B��`
�])q�0��8*��ؓO]����4��0�.���W65�\%Q�!K�H���O����c�,��ӷo��.�yFp����^��G(%�ǽ/���OHl����Cse���Y�c ��6������EWϜ�� �L"�Iӟ�� �B���  | ���U�!�ll�AlDP2ڒ�'�0}фq�$爨� ��Fi/k���c
���b�Gi��V|-��-5�[c&�ÕD��U��`���Q]���̕xmdgI�m^�wlqk<�1*G�m+`j�N�л�~iw�}�aS�c����Vҟ�h3�Sd#-8o�?{6
�AC �R�M�wN
?#��؅}"jv�A�rz�_���F&��g�k�1R�W>r�E�B+�E�Nwg����F oP�Z�JȤyYK1�X6����d?1	��?�Er�X�_��9Y�>�1n~`e��d��	��G�J��q��ֱ���[��E�n�b.��ۥE��s!��O���ֹ��]��2�]+ϳ+���4���8f!Q#���8ffi���	ԣ��A���~�ڪ��FH���Ξ��A�{�Q�1]�L��r��)�e93��.˱��﹇0����W������2M9��)��.{�mN`���hv��[�Ƿ��S��.�LΦ7���eN�d ��9�SǱ(�{J��J�qi�
؋���<$@T�f�c�G�jg������5��7�TF�C#od6�l�	Su )6����~�8wKB@��wz*�l>�yL>��x�kУB���   � ��u�!�,�U&txH&�Ñz� }x�Φ��&jf^%���(h%�8D��J�y��k�n��$�(��f��O�@�D�@�G'��jrɀ5��?�X�,T��ėA� �Vٷ�S�/�I�6�>l6	��iݼ:nˏI'�pGs1�	W��s���ݽ&��F�*���B�"�ƣ�r��A�Vjx��'��X&�G��;L��U$�=�g��f��w鷿 C v�+���3u��;�'׎��v������0���@`PS&_����i(�w�g�|���D{=$�\�p>�<1i�����2��sXʩ0 m��#�rЯ0+�����hhd�d	��p����D��5�d�w�T�/�q���)�hh8��M�,q^��CE���J�3JV��k�3p;9��]~�Gd�!I�	�m�0��顺0�/=L�04�AN-��ww�z��/�^�w�?�M|��n*J����ՃBq�ެ�O�ǔ�M�C���,gW8�-T�&b>���Qau	�$���ŧ�'������G�K,��ELʣU�y��s��[�����%�_Ѳn�Y1�K_�%��eT��c��#M��$|kB&F�\I��t�n��# x�t�0�ls8i���H�f<�s��.g*wC [  �%����أB+�O   # �B-�����zH��NN 2�h�
���xD�qDqO'dB�X'�	�Eia��H��v�'rT��Y>T���"d-~�&T@֙+*K���rND^q>2?@��:~Mtf��. �����_�.S�nw[���؊�����hQ���6t��c��,x����@�b��ϸCjۤ��榯Su�i5�Js��lǌd�-ƍ����rzrP�԰޵a���`�pi��:^P.���=a67M�Lk»������Ў��^s��	L7Ba��E1�rQ���F��{�Z�.���e?Kj9q�����p�=�i~�t�"PՒ�����,hm�ی�ȡ 4�M{f(�� M	F�J�9U�Z�E�]^>2�0�<�������Η����H��s8(�����=R��z��+�����N�!b����y����wYQ����G���ӡ�04���C�O��?y�6Aܮ���o@��K#�%���� ���h����_n�rK���^�� :�ܫu-g,MDD������%%�f鐡aѮ��`�����I] �E~����������!���D0PbDv�` ^p=�_�;�KG ��Q��C}=_Et�A���?�H�{6K�s �v�����hh��E��Q}n�i�KƹA^J��A[Z��i,�/Ӷ0Bh�D�XSNDXJ���c橱8| ��>�u���$���\���֝ӡ���nv8      �!����C��.F��!�A[��Iv���Ң����V�T��/y��#�[�
��߻�x!4��܅�;hM�Խ���5�/��SWL����Ȗ�kd� ���<�g��KP�`��ɅO)���3�;a � c��o!؀G6c�M1۫s�����U��    !��"�D�(�"+�L� �A@2놔Pl���:K��9@]�e����"Q�2����\�g��<� q�M�`a�rh(���!(�N8������ �t>�����o������
�B�p��q7�a4���!�c/�"� &���\ �~�)V?�����2f�f 0  �!���İ� ((��� , �V����g ���x[����d+���o$c迡L�AT�e3hΤ#��.�S��}��8&uB�\B۬�]E�d��s��@f�D������/`@��[���M~��.%eBk��\7�	�(X�
Z ��}<�K��B���쳕w��  !��ƃ���0SR�P -D�Q��T�Q��ry' �F����u��o�䟅U ���HJ��$�2�f|��2�s�:U7��jYV���!,]o�����'�J��,��|����[&¡�d�Txt[���6P�@��!O��)7�n�Y2V�~k�}��ߋ�l�    p!���ñ0�JQ:��#  ʕ��_�|�-zD�ϖ�X�Y��{�1C�'P����^b�?�~�����W;�q��X7�1��p�6{��c�{�P59��?�*�2�s��tB�>\紎���e$���.��0� ?:7��3}Rޞs��o矾s��     p!����1hq U�Z�h�q��
#+��������tє,8%��?�i�3c)�/��������lB�,����؉^�J�PETLM^m���pjt^��0
�UIAsL~��<�#���F|U,
���o7��e/�t���$!�A#@��eOJv��x���g��uy^( �!���Ab0�a~K `m�t��+&%��Ƿ
��>��˭�Q�ܐ��>�	})3��}K�0q�%L��R$+�/>8V�]�,z@��U>�f�88�V�O��-h]�L��-�=��A�"���{Z�O��F�O�H�6�:B  ��OW\�;��C^%�}F��T aA�H^R��n�  �Mā	J   �������C��5��/�ώ=��E�`�`L6 '���lF��#@�|g�1Y�F�\1��%'�N��k &�^ G�������q__2�:&�]���a��£�I���Sҟ�� ]�"�{�����=��W���#�l��W���n�4��A�}9�L�5�~~�3��̆l���2W
Xsq�i��� �c!���}9���9ғ�T��\� �'�#
j+��R��s7�%�	>�E�Ԁ�!3#M������ շW���5�L�@��'R�Y巀 �����r�m�w�\�����4L�<�ᛴ��~j�u=N}�!:��;Ыy�p�e�ag@��af �p����k'��x�	JzE5߾�Џ��]\3R���h�2�-Y���˽�k>�t�G!b�7�%����\��M�۹&�hȢ.ro�xtjv�q%E��k{8C7vě����a7D��ϲy.�L2d.t�*>S�_���~���}��G��E�/��&�Z���lU��IRB��e�>0�١XSy�8��pȊ�H�"Jj��jjZ5�@(_��Q�G����Ѫ���~��d.·;�$Ȭ킖�b��DT��}���m ��F�rqi�@�l}� ���B��<�Z�7�+��L��Ѽ�{64����:�����aV�=����-�L@:_��͘����`OR��;X��J��U\)�d�W�SW뿠��@^�e�\��i���3)x䍍.3�q�`{��Yzi��r�hn��kc�4v�+s�OS�F�e���c�"�DG���\R)��峖�s���#-Rc�{+y�dmj^��'l�����g��-���c���C�Q������EuG㕢~�9�����I�]����?$%���ӑt:�М�G��""fd���6��3�L���Q�F]���Q0�����P]r�m2�^oG�H�],�r"���w?`����3f�#E����؇�� ֮�<��>	�p&�$m�C�Z�cB�2x��Z;I�?$m}Fc^>�x��i��,7�HofI�����i��ϼ�!�?42�	<�*�^7��徥tN�L����ӭ����������m\͟[ޕ�����#r��m�f�}��1��%�!*\.n��^a���Q@�7��3�s��a��Exӫp�[�Rߎ#/��s�Zi\�XM���`q�5V[z��ጼ�V�b�?�Yd�"���8Rh��A��֖�Wg<S�z�n$�18\X�k��_z:����E�l1����V�ZUx#���)����e�x+�Nw��!`���Yx��ʔL_~��J�hs����}��M@��f�p?X���
��(������/2������b@o㢘�����~�]t�{i@8G4��ޫBl#�q�
JEn��%��8��mt��=��Ba'�U}\��O�k��}sS��쵠䋦��|���$�U6-e\ܧk���j��i��i����A6\ԉy�>�&�7��'�7���9�m��-E��E��)��Yjn6GZ��x���'��P��`�zKnk�\�=
�˳+��QUu�NT�>����c�-��L!M����oJ��{8�&,Le�~;��I�2�+�۽jJƃ���U��ˬ��=��Q9�Xda༩�����	�� �Y"�N��#;2|I.% h˥`���j�w�^}]�-�F�L�{�5^n���t�� W9f�UVB�ȓv��<�+Ts�|y4���B�uPL��&I�)��6^^j�l'�3����
N9�\��R\���I��@ƴ!�5��z*d�j*Z�:1��64��,��c �@���H_}��S��}-_p"����nqp"��	��U���?������
����'#�,�U̗���Ħ�Y�� =JBZ�˚��H����2c�8�{��x �6�����<�r�xU�)�X�H����f���5bΐ뿯��Gf��#�+͌��nE�fI��S���*�l�1Q�P�� bj�������
0p�\���>����:��xX*�Doಌ�_n%����#��,fpxdG��]?�6�Pm%PM�I�#ـ��9�T�T�M�E2TT.���Muo˛��U��h�6ӌ� ��>)%��Ɗ�~8���2��
Ϙ0ċד1��4�`�ǻ���[/ͫ�+�%��Zk{��N�}Җ|c�Kd�n��*"��+z\3�S8����q��g�6��#k�[^��E����H��|,s�������0$�K[��*�q〷�ue���QJ�K�"��2�3�9��ذު���А�	�hN��ǰ�]щ��+� l�����ԅ܉���v�aX`_���a	�Q��x(�b��<�#�-�P�aj=��Ϗ�^������/�Lz�0� �I�ۛ.ؽ_�[_B~X�D�8���N��i_��j'~�B`�RL��؎�&�@r�i��n�l��L{gAb�*-�{�*̕u������wL��H4��D� D��1M�B�+Ð��$=��E�fn���Q�{y#�u��}�\7�����Ӂ�w��>�3���.�^�By�!��~I�H�(�L��Ι4Ф���q_Lc��Qm{�F�0�#G��>W�i�Z��e�D�����iO�(����Q6"H�;e�i�wF�#~�V_|[�F+qz�]�]#9��/	 -��)�K_j�N�/���{!�]9�X�|q�2g��iz��f��B�qu�������I�3#�sE[g�^��o���N�/H�N��(WL�ҵ�?��h��.��H�B�=�A(.��U3\v
��kt�@G�X�u�-{���1�bNRBh���1a��WY�H��z��]�^��IMCš�ʜQG7�v�F>�m�uH���y��:&�,��]y�9P8�"�p���3�Y.�ȁ7��WOGc &&R0�p2�s>���]/����.b�}C�E�>����VflP.�.�f"F�!ZZӹn���'�� r�#�|Ka�vww�c}KLlL��nZWм�Ge�5MI��֭��J�"Z,U��jO{yL���44I��mJG-�D|�M
g+�[�IX�*2~��-��7^���������2��Q��±<?�8�_BofDl�r:�ܬ���<J��us��GT�[�}�z9�J�نb;v!�C�I��&�~;�U������.5x�6�m�XĻ��<�������dg���5���I�N+hԉ�Ք�l�F�|�G�$�2����H�5��B*��]�<��gK��;ߞ��E'~vw�ꝕȜ6����ۮ����f)o>˶��?�>N1̓��Wl������<,�ΜV��X��k�y��\gl��_D�۶.�����kG�5l%8�� �>j��v��������#����h�>�z�S؛oޚ��������u⢶�Z��?��We�?3ww����d^сU�U�I�k�d�k���k�9���ŗ��N��i���_���/�����?k}y&���}G��	c�nt�DJ��  B��'R��c�:-$�xJ#��@����ٷ���ab�_��
�_��Sg����{ 44!�N���R��
�ϣ����,Rp��{0���Mx�I���V�C��������X�c���wSQ&�=3iyczv�F�6�s{#z���SC�W���a\�K'-u�ҕ׍?���h9o�� �r����"E��j���I�
���Nq3�H��_������Ġ"y�Q��03�w�,X�a���b�r���j팤v��拪ZrUȇ���E�t�
ډ �z d��5z#��_�=�m>��*mZ������{�&�@Bd�A�5(n$���`ʻ�*�v~P���o���X�gEUwC
�: �*"��pᡭ,j���h�}8�/��v��7��f�L�)�s֢7R�w?%�?T��e��v2��T=`]������G��ˉ�;:��[7[$NC�$P]B;�7o�n���stw��I�^�z�Exb�+w�?*J
�F���wJ7�M��`����M���_*�4y��sb�)�|��� ���InY���U;>��ȐQ`�K=�.5:���ö��^�2V�V����g�pG\J��	m��UH�owɆ�ء��Ԍ���
�m�����	6��ʅ�/{�в���,�Yܔ��)�Vng(dI-�
��a�
|���@=
����$���{WL���^�y��j	H�ͩ��'5�RtQuAU��,���c�s��@�3>�8-�/��Mj�
��Z0-2`ҕb%턳��� �H��*e����2k���Η��l�N[�٫KNKZ���<0�+n\��;�{�B�L��ŢV�����4�Go �H���k3]x��^=��"����ُUu1{�ʋ��J�>����3P@�[+���	�`3Z��ehx1��Z�ɔ*\�Z�|ڟyᰘ��f���f_U7^9�n�1̏#���W�P 6���� "�t�ޕ����ZBuf}�"�	��\�����ӽ/���%H�؃�rԖ*j�idx�$�3�FZ޺±P|�� &�#w�#�i�{���<�
�}ӡ��1���z �!�k�Bہ�  � ���U�!�،�"E��\@2��� (�E�i �������Y������c����=��c�Vso��Q
��5 h2��Ę|���r�}P1�;����\;+�a���[�!'ٓ��ur=A!<4m	�0���Z�M�H�"m����߇L�e�3��y0^@���8
P����=Zn�~f�(H����Zg{9�v�o�l�[���D�L�ׂ��s_6ʈF}��#���
 �Y��AS,E�#(���|BS�zF��{¤غT����1>�,|��{P���g��I: esFi�w��s`� ��������������h