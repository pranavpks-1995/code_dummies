��K��s5�F�!6J���TJ�e��ا���A	|� ��c�������O�U���h&9��������o�wt�tt��=�(���4|�7�uYϬ�2�2�R��b��D��r�>o����ߕ�R�2lI3;�N~.U�^��u׭ne
��!/�;�����E�\���!�8���7�m�CO)�D��d�A~Cec@�G�dÎ���Y��}s۫��tz= �g~k���r�=?5�~$��8$�۲�%���z�r�hD�*�(��b���� �݁q�.qk�ʨ��zL���`�7���۷�D���O~nB>��㴶�2��X�ֽ�d���c��k�w���s���5����rs�1cOFJvYߊ�>+J�F��4\��>b-j ye��X���c
^b��F�u0-LDZu�'�?گ{�\���$�#�e� �g�Eoݫ��]������������!����{5'��g�3>��w�X|��;��	�$$]�����]h�8�X�h3 ������ؙr�	�������lߗ'Æȭ×� ��eV��="��||�!���ޭл_��J�1�'-��%�T7?�,�o�5>uA��]��7�0E�<��Rn`E��k51�as���	;x�SV���2^��arwWZ�u �����n�_ޝ\?|LG[�����,�R���H�R��K�
30)mg��s��b�p��l��9�(�|`�f"�)@��ۦ7�۟ז��^ȉT�����'��?�y�����?����U��]�g�Qc6����������;�D&xi,PH���e.��!��ky�P$ �I��{|�9ѵ�
i,6�ɽ��ă"�h��n�s���K�嬒[.]��$,�(��y?xk�s�)�3�,�J��q��1�4�^��t����!��ݨ�����}.s�?1�8�JV�����eG�[����1��/��]����'�`����s-c�:^��J*�lDb& k(���% �����ҭo��5����	���-���2r[�×m��]zۂ�hc{Q��~�R�� �;����ȮX������*�^��!���-�������7͈+��Q��� j�Y,rZx�j�JVd�m#eߤ�$���eH�Ye/p2䞌������M��rO�2��[��rZ&�0/6�%��j+Z�{Ji���1�ݐ�����:��_��Zn|�Q�l)Bk�;(�p�������1��C��⛩�n�����i�iB��M�l%rN2�	e��.67���1�\�b%T^(��ӌn���� Y�&���o@N5�Mj��˹xJX�n�F:�k��*�����g�n������.d�Q2'߿[��%���B4Q�igt-IZ�>*>�lTfcAc"�����=��3O��v��q��F�)�m�d���.
�i��B��oZ5��VEv�
������ a���痟����rQ�;h�='$�N���wN߁���V�x_f�xW�����fh,�z
n#��3����-��&.a1��TX��V���x~\K-�6�>$9Bq���=Y�Y�sg����bd��iC�����˩���p��Ikx�]g�����[�
ê�x��{ s��<��>�X�<�wTq2&@R'�!;v�����f�rk�A%_��r+jW���(ː��>9�z�}5AA�c�+�3���7�:U�J qL�� ���$���}����m��N�\�;�.uv����7����fxk���P]]Ѵ��yE�۽�H��}�7���9"c������ٸ����q#7&^�^���&%��*�`�X2����-�e�x��2L�ç����L�*(��u]�懽�ĉ�&�VgRc�"+Y�S��$H ��J#���g�@>Ʊ��:��&��\`�[~�TT�a[W�W��k|af� Y �ݩ��\M�e:F�!��-��S����� Q�����Ӛ.��������4cJ`ի;����7�X��'N�jl��PI��P(���mV� �ϻQ2s���|�{f���v�� ���<��p$@�YL�r�V��d�`�% 5��������"{sR4,y$����\n�t-���b��9	������Q�����gf��0�{�`QiVM��K��-F&q� ��'���������3��1��N)t�ǳ�-֘�}�@s�ػS���ƶ5�+���Y����[K���}�g���^
����ݭ3��V�Z���maG�6~"�fR�z�D��P����X�͔ � &JU�.{���C��|�ʺ<���,m �ˆ%����F��v��{ :8�#� �8Q1@C��&_������5�=O�,��,0O>�RM���Bo�X�`�A�ު����Tl�dIi5��Y�I�H�Y�М�ө��`?���D��  � �����,t`���.��b��$�ר��A��V��F]�-�͊�}�:�22��[�����q�N��k;�p=���8 i^9r��,����ɀBb�o��v�ʾK�����??׭9f=%z�mQ���B�o���i�P|����?JrM���d!o#;s*����v9�����K~6�R���!�K!��o;eմg9ʖԞ?N���8D�SUSp�a���S�O�9��*��uo���V.���0j�K{�G��ۡGt�Ae�����G	d�S�u@b댱�j`�6�8TY��tl&�k��G��@7���̦"+~���$t��>����F�s=��0<�����n1�T�ͭΩEs�*$�Pj4��bއc�;�V�{0s��aA���J֤0鍺��'�i_�_�����@�x&�D�h���p�����Im�����u0۲}aדe�U6|�al*�8��>m��9�n��e6e������)�-����j��9R�	Y_��S���"������ZH�L<2���l5�Ղ��0;����e�-���Ԡ�����ȕF�|dz���a��F�/�����z�3�����Ĕ3����Ai�TӖs3Dɿŗ��Rj*p�l�ik�ߒW˪%�/ ��E����1�}&"I����u�W��J�tK,�:�+F�:���B±�C��i��)nO��Z���}<!cP����k,���a�Ǖ� ��N'�G�I��U��9�wA�;Li�K��Bv%'��U��`���-"h8fq t�hjH��m�NQ/��^(�#��y�J�,�Y��ÛE�}5��h�mZ�q�Ȕ�Xy#��gN
w�֖��� T�r^�7�҈9���&�6��#��{�j��"�L�z��`w�������G�:د0�wk��>����9D�~"���Re+X�6�Ml�>�,��#�Uq���\�A/6����6E�	��o3'��4��\Л�C/��b�d���ü���� ��Z��RL�*l�oM�G��X�G����=����
�h������� *{�0�*�#]M�����<��#��Do$�����Z��P� ��8������m��*�tc5>�1u�h������ӫ�8貀��]2�y����P��!i$7.�@3�)��/r�Y��7˸��E�[    �"-W���+��Y�Y���@8"��^b?��f�����(*��l�~�l<x��ć�ɏf�	=����Vյ���"�Dx��bI*no�A�`���46�┵BXzx�mx���jA�.�t)����,b$*%�>�J|K6<Ӌ��2|<�y�K�����B��;$�^<�yt��jϣ����SD�qi� ���4��UW�U+8�k@cx�c7���J�D�H�Zl�]���p�(o����g@#��o^Q���.|r�Aj)ި���&l�<�������:[}r�T�7`��1^x]`	�,G�e%�?�d���-�C��D�/v0���p���_��٢q�F�� ���y\^ r0]�%��.�G��x+���)��T�~�����;'ph��|��0��=����)Y��d�WK�5�=
���E!�[���!���V3B���hwtǖg@ы�{�(k����!}k�Ά����m��Q�@�q;��le��3+4� ��w&����%��� ��WD��_]WhqL��>7�.��wfl�����p��@^h9�~�Y��7Gb��gB9a��\!��JS��kW��y=�*�K���D]�[!5��HH̵�#i� ���J�zAD=��^��m0]��e��d�?�X������:�&�R��+׷/���MW��"œ��tZB��x,e�����Э�F���}�:�k�d���߄HkV���k�$�+%�Zjv����b�����>���t����	U�Z	TN��1�j-ַ4S~�q�	�~g�i�I0�?����v�%�f����R(7kio�Q�B�G#w��%�r1oT��)��v3^�0��$$܇�u	��P�U_�\J�+�o��Q6Q��^k��{:��Yr�Qs������R'�Z4Lf��l�RGGf$cؐ7����Pڬ0��ڰ��Ü�`�&!�Ҏ�!�p�G�{3΄Jg���}5@�����ns�i����uk&���5A�a��"    3����^�i����ǏD9�Bg�O@|e�oQ:�:{7Kt?�'�?��݈t��!�3�A���X>8�ho�� *��#�&���'R����R1b��c�8������Iܕ��2�L����Cm�|�IN�B^J:�|�z-������Mk���&a��<�{W��fk,��*���������h�Sf}��D�eՋE�5\�yB���tdO��P�!U�_��7����lz��B7o��CER�g<T��´�W6�� PDF��1�  �� ѧ��EZ���ᕞ����!K�F�j��4��UWWE[�аv,�)~-�)��+J��,F�n0iea��j"�&{�ys��
���/�v��*':��|m*r�8�F���z�	�s/@�r�#f~�^��5�?`�(�����!�dop��β��CԮ�*�_}�bI�;LE��l��y:\]���!;����ф��D�dAҠ�e 4��
�>0,P��\��JЧL��T��-P  �!y���±A�pn�d�Y��Z�+�=�10�v���~W*�KK�����b�b����PZD�̳,��r�	l�  ���-] ���\d�����j5�#U����A������pY�`XJB '@�X-����A�
Ŷ��]����iP   p!��T0�h2�Ha@(����Պ}��F�Ց���c,����,��p��� ���r�]�O�^3M������g���P ��oKH�'H��,�D���?B��]?>���#uHR�~aiL:B�����b�����vF�c��}� 0   0�!)���C�l1R�
,h�@�ZN}��������0�g����戼fb�z����1����@j�	6���K�%S�	�*���C0�b�&1�WG��aK��j`�nm.�I�~�B�Lb�Z���А>0�ӼH��;�v?}�9��Ҁ    !K�KZfz�G�.m�!D@��b̺]���
5�YeE���&���wv嶍�L{f8	a�ùK8<�i4���5;��R���5B�"��h�S4������D�r���"=���ᶁ,oxVD���,�r�L4$��s�0��<pm�92M+��}1+��a�G�"0���x��e�HA�Ho�r�0 !y�)�ı �&�*FX�n �B�F��6Ȋ�����0�j k���#�����`M͇@� l۾��oP(�  4۩�"��.W�����q�mHZ����Z$F/���%��3����?�����}���:"�{t��7�=�s4�   8!���#��``R�Y,ġ��5�(�@'�e����FLn�
����q�A���k�����9%�b���0A�%�)g����%j[��������d\�xȋ	1�M��	*��+L�Ϗ'�Z'9C�y�p��a
$�	�Y�!TO}M�Q  !���`�L�5RC`7� 7=΂C���H�D�1�%����꬜Y��9�a\0�ZH^�d(+��B� ��<��D�>R��Ic@��*���>rZ$�o�#J�c`Z�7u��9Q�wO_ۮ֐ؘ>Ό;�4""������0�ϑ�߯�ך�D 8�e�,   %�Ѱ�UW�C���jn�����$�hXD�‒;��;���𦒚O#��ǃ�Pf�ʸ��i2��2�[��QP�3Z��7FG[3O�Wk��,I	%�Fc鱞�ҝ��Ƭ*��F�Zګ.�iH�=�s��M���h�gj|B�L�{e7̱��?p-܇t����"B(#��!�z/0�o���h���Z����8	`���M�im�X���\k!贁B�3yO�)����%W��ZB4���B'Qak.a�Hj�g��{�A���36�'�<����s�r{8T3�� Ô�1�(���[����,�'҇N�>���+L���iW���������оةtl��R?�R�L���~f�eLr�)�Ƶ#kne���~�q���L������9Q��)A��B͌�cd��
Ė�2

�H�Q�C�޵�jL;/��F��s]E���������4��O���Q�~��,�|��Q���F�q`U#�l0&FL;�r'@�\�R��F�Jc��f�~��x���rԵ���VO�����W�'�:��N�`��l��̇Vl�swRS�J��-��	zwNg��,	wM�Έ��jC2�"��sJ�ǶZ����`�gy���b��m�NVHo���DMz_���rǝqv�4~쌚o0�*Q��0І��	Y�vW��24Q����/�J&��e� ��/pȀ���m�Wf��ܸ�����6��~pּN�L��#& �/�[	��eN�H��5���t�����}R�5�bf�#sT�P���O�C�0�p����!����_��rt�.����&�޶�:,QW�ƙ)0����o<�b&Z�Gn
�hs32�9��f�5IDX3�o����΢y���@��nj��ԂNu��>+����jl���޽��T*���9<uEa��U����u����n�m��T�C�|�SZӿY �O����Tp	��t��N��}�N�Jܲ�]V@�Y��(d�D:���P^���:P����PrӾS'���Р'͓�d�{1F)���Ĥ��o ����w�XEh��*��Y3���X�M�>[�kilS>9@��ml�S)�N�u	�T[�I��p��*���S��(g��TvH�,�"��3�p�����Q.\���e6��$�a�XT����������8Ok�4c9���F���yR��'#x7��,P�	Ħ\���q+8� ��]�O4����ߧ�GЎ׽r�6�+k4Yӳ��u���f�[�k^� Ơ�PjKF%��؃���(aW�[�i��kMd�
C9�]��g�Wr��}�j�-Om�b���(��V5�ڴ��Iz���s��*���e�e[��
��/�i2Ha��lL	���it=O��#���-�@����ˈyE���NWis�^�A�d�DV�b��[*-��5bn6t�Tׄ�i(&Ayj~���������N@���l,���o�.��|��u��C��}O�EB�b���q]��a"0��-D,_�3U.�U`ɿ�ÿ�o�TQ��f��7�,\i����=���rۂ�br���	;,�E�FKh�WD��ot�����>��O+>f׽W�M�GP_�v�, �p���o��8���`y�y)��2L�)�(yϯ�2B!�������z$f1�	�IX8����uP|� @� �1ai"�*C00�nTG���K�7�@!��~����'� �?�˘��������K����3[^��q 5��W�,������Qm�f)x�A�#��!�{xrvA�5�X5����z�>$�>$��A�T��<vf��F@��b#4#�׼���$]���yi�9�}ʫ�ۤ�����$5G���ǥ.>���\=Ut��Zok����?}��Μ��?�<�'�� �*]��cz���9֥�^39�W�xV�{��ɥS,˗�5>��8��nD���W�/��s��	��D�56�^ˑ�,�J�z�o_��i
B��i̳{L�J��N�E�l <�ȉZ�|l�Y�����*�j�=GQƼ�~������!T��ئY��� ���+��&�|V�U��0���c�hN�>�A�6�`��>�#VʎQo��Ӥ	��G��E��"�:y�PN�w�,��5Ҫ�$`�U�ډ1���D#�<�<��xа�x��y�W���:�@fddu����v������ߑ��Y/�b�%N��o���0�\���P9�
ĝ�k�p:q�}�j��cKFz���Ѿx���)�v$?^�������b������{=|U���,��E����O�zCo���@�?��ٳ��kZ<�b*f;�"�J˿���<�����W�W{J��Z4��L���z�c'���I{��B�5+��=t.�˻k-����z�.�<Dq1���E-?���fP�(�L 2#,%�ހ��=����P5ma�g??0�'ۚ����b����@��Sr֐���C/���3bʠ��9�D��j�bZd�R��-��c�Ά;:���kw�����o��fř�;R���?���G��%z�U��H�G��Dy%�&�.%Ӈ�)�)�;�)o�{�p��� +�|pfg��,�<�ӢtB��9��~��S	JfL��46���G���7�3���q��XF����U� �%�r��QD-� �m�v�w|K�A�s��m�:D֎�w�@˝�S�᮳��q�|�P�JE$~�7P��5-)�S��?��45�3,�K��01����w���ج�1��ŚM)�o���\��?e��ln,�)ز9`G�
�V���d.�����-�;b�8�BI�ç�,'�G�U.�a���Ղ��*GWVX��>v��2,n��q7�o�^B�hn�6x�jvho�X���~�/�E�B*�m�p�-�)���3��΢�%��~6����3^�*]���P ��5^�jF���6�|�l|�ў]�%)	��Ȓ�W��]r>曣�3� �|�6R��Z�*/�dx9��x�D��m�pʃ�aG ��k4s������R߬׿8[G�:�o}�Hk�P'�� W!�r�F� ���h�`��M�����М!�3�84o���h[iZ_\�:8�䬚O�~C�)�:dD��"�.�����i$e#�?��&�l��JrV�I+����(V!�۟R���3�0#�h��%QՊXͯ�=ՙTo7^�y}ɔ�ɭ��]�6�Y.z�ܭ:��T���%?��;��(�J�V�]P�}�_[<�@O��z}�J�o킲�^��E��W|hFi�i���z� ��ZPTN'ըJ�f�'m<��'0�TC&(|DtZ����]�?�x��4����.������˙����"U��\�߄6��&q��E�)mo�
�n�vp�T�r������b����4
�Q��<����Ia��2�'@�}�"�K����G��<����