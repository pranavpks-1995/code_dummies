�I��5�N��!L�@�Iڂ������S��iC��^Tu�(�h��f8��KB�*߹O|��"�Q�ȋ���I�#L̀q���)�uK��q7��Wp���Zfn�C�����|��M�n1��]'�	�d߽�����N� ,�������0�W�T�~�c�����_��*��I�FQ|�M�����	rF���b�.�𬮵-�D?�#�P����1/rr��ȱ*إ�$!F�֋:��O��,�#L���B!!�݄R�G,ÞG��!9��*,�Q�k6��Fĵ�%SW�:�LM�\y�@E�������=�?��5��䝝/����`����z�G��oC�m�-���I�S�*.�e���Ӯe�=�sIu�j��s8�d�x���!���T�<�T���Y�ASEW"h�>8�������2��$����Y�>tKL����tK�4K�]R�t���?������	_T��W��f����N2��� �
��dK�����Lvb���%�8%*�>�{����1é��&f�s�!ة��ӚLe�����)��h����*��=)קa }I"A�Gݐu:�o�*:H�Z�i�b�Q���x�t0��v���4��U8�]�Ƭz?�'%;��4�#� �������k�AX��sߤ�͚s��)��&�U*ip_��A����;IؖPwg�|� �fն��g��aX�]���OCC�>�=�E}R�m�����ک�D��`@(jG�@*���Lk
�@"�'~\���	ˁ��d#G�-Lс�"d�L߄�)�>ڨ'�]����y%%��J��/�$b�"�OO�Ҡ*�EUp������V�~EZ��[8�;��a\	��_	��y��N�#��s\?ׁL�d�R�J��b=�;�n	��Rn�H�"H��W�Ö78=jT�	���\^����ԠtBN����Q�B����C0����0V"R�*C�Q�[�t�6(U��%5�Z�tF���i������7�Ķ��{��`yP"��8�k��zow����ͫ���Vmy��q����3������?��A!�z�#�?�2���7��}9N�A���(��dɡo�0�6�R:nnX��N���$����ٹ�8[Ӯ���$��r^й))������V���{�V�[}���)j��R:jp����u���d� ��K��l�����D=��e�'�Ȓ;`��l��s�3����Ct
nt�9��_p��AGW0͒)l#hۥ�M�x�� ���՜i#���:�肖zuߡ���y�h�C�����)��AP\s��2E��2�:�P�ۀݜRmP:z��#��C�/�|��D�D��W}�h;cV��)����'HVc j�rеd�����z��F��h�n4����
�S�Z���TUj�A�`�����~�`��@=�78�(�fM��)�#Ij�>�S��vh� ����☄�XZ���F�O�*��� �dt��e���wś���s���J��H��7��A�t�(������}��k�]a�:'Sv�!�P�������S���B�`K����\p��Q�w�X��(�<�X��R���.���魜1�>� lQ� ��3�MB#