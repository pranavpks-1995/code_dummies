�o�x�3Ȥ2?���e�/����SV!Ip�ϗ� +`0��8���_��H�1�2�O�J`[���0��ۦ�0�,�p5W�eg�[���h�"V����,B�7��
�[}v߂��`  p!���,�����tX�
����ܗ�9������:�` �b&P�<�Ϭ�
�s�9�?O)-��z`g�~���a�9�D�C��@>I�����3q�Kό�����1���;�����B_�X����$�*V�r������>P'�HYL�#  !�������Ĩ!��mR�R�����c�i��1dWlN0c�}k�N�T�����s��w��= w�ɉK#E`<3���:�2�8tڝ�[k0A����2��O�X_/���1�
MF(>���Z�E��-��Ƈ^�*dB0Sv������8���  !�ʶ* �|��i��]ĭ8��ϰ���7��`;��ߖ��:>�F����˂���j���c�U]�}|T�{^}
�7����
)q�-b��u$;�$Q ����>�h 0���f������B��霹}s�  !�ʮ�a	T@F�P2�d%K���IuVcO���м�5�������9������RW�mٛ	L��/����g��^�Bn�n�m�6���TK{��ӌ�q´�{��O��(�q.�EE���uu:��\�E̗���:B�����s��> 4 !��"���b�NGqx�V�.u��R�R~�L���B�N�F�7��&����4f�ƒC���4Y�jI��M֦FZ޼L߳��΢�i��8��s����S���҈c���`��l>���  �J��	a|�ƴ��˅$H��  p�S��y   ~�8����C��\��3�������4�G����~#2$�������qB�B2�P�P)���G~���3�+��e!���d�̎����A�-u�\s�]�+���v�y�4���.��_N�ɶƝ1��!���~�zV�T�S��9�-�J�;^���/nmJ	��1��m�#���
����+;�B���T1��}��	D �N���0�����p΂X=D�:����?�wf~���[)>B�?�