�ڭt��?(�x�92o��l���*���I���5�;�4i������ĒK����oG������s���=j*B0�{`���b�O@����ھ�x�w�W
�p��?��'=>4�SV6>Hn����l{��}6��}�K�^��穋y���B�=c
d�\�d}�! �^�ܛ]��߶���� � ��/�m��
���r��fE�C���dm��;�q����ߡ�X�s�<�I����#����ݡ �.S�'���y+`'�,�$Ò��s�_�M�2�8������~�an<2:���!9n��hvV�zsa�B��$;��J�(�����"��1K`"i]'VDO�;R�W�η�������c����]n�=̒���yI��ęJ�'p�3u9,{py�,{��������o���|�O$ݝ�ese���9VD�]�ڄS,��H.Ԇ\+��-�(�w4~���?����o�7K���s�%\�L�� )zy�{���ۏN�!�t@��' 2Q��2�6n6n��[�
�f|���js��$�����*���w4���)��[����>��y�lbRE��eq���� ܋R���dsxoQ�-|�d���$W��3���D�G�. q�z�^.����F	-�$*L��fK��`����$P���v2x�$�/1M4T:��=[���w���_[_�b���#:�|-iX�/�0�T�Pn�r?& -�x ��!cd,���s7��J��@)�F��+(Ί,I����7�`�������4�e9�e�|������=�z`�W�$g�f�1f����C��  ��'R��c�
�60H�@��