M��0�g��-���rL���,Ь"&��y�:e����e�HN���	'���#E����1��0N敤�E4��i��k�;"yX����ɫ�Bf�AY����*D3����͕��o:f�_6V�?+�j��+��r8M�O'Z�R���b�O�x��z�m{�\�6,������v�v)��ݪk:AȒ�^�;���`�^&���>���lG��g���4��M�6���� %�LRLc}H�bH ��xl��C՘`@�r��Gzst���s��v�(���Ap��hcRZ(=a��n�l��y�P��E� �    �f��F:0H
L�DZ��_��(� -� }H揙�P,���=*�:xHMZ�pui��u� g!��Dq��s�(d�擹��z��a�.<i������+���::oh�0d�{��
`�h�ʕܿ�!�	3ʊ=~w�u�nAݷ�Q-Ċ%v��]�RqM�م&k��{)Z� �Z
�)�<��a[4�?�7 KA��n�6Pg-��:�ՐD�&��!���Qfq���	���5��G�p{Cp���6ҬK�"/_�P�ƹl�f�����χ�?��L,v�����4'M�g@�z��ݧ�_wn��P�KƑM6w@�
����S����k(A�,��'�����T�C�m,�Z'z����~���7��C[8#:�s(4~�f�1���p�&��m��+��j��cih�,ì̷l;P�|���r8�J�v��N�����kL���8		F�`��>�JX��6�\|��讛x��i���-V�C'�ݧ^ףM5mh?}^\@0��_���a��t�[��'M��U|68F��0(w�6�?��rC8/��۵�`�ʙ�5\�9��U�_�:� u��NM��YD�-�.9��-� R�Qq_�x���e��:��6���������f�~m�*���>��|7��~��9�ۓI�B���\�E�;���7���:?�,����4Ì��)�}	~T�Н�,�%_@���XhS�N��/M�Gk+�F<��9g��J���$� �L?EB�^GRh|K��^,��DQ�Z���Ob���A����$�_惹K�Y�������<Œ- kW��{Un���e�(m2����}|ү빩b����x���m\M�ֶ)�4h��t�{�~˱j[*ܳ��e=�@=��Ӕ��S�{���ot��	#k�'�p<*?5&tD[��j�&�h�ժ�����"ik���,�gF���4K��3�K��!��q@�eфp�_�(l���Y��5C�8� ��O1��Cd� ��Cv2���Ln2	c�W����2�=]i�{���gߺ�����#������^7X�>hE�hBr3b4���Bb0x�_�y�N�7p/�
����)��C��}���2h�[CK5 b[�)0;��34%C��1D9Z"3��rA_Ζ��:ܤ>rP0�h�F[�Rb�5�c'#-�>�Hw��k&��?�[��M�,���%��5U��[������:��nmbb/�n�A��G�y���hB:����7:��ܣ6u8m���&��4V�/��M�\fd��Ҥ��ݷ���E��f���Ǳ���!�J*�.���"4 �����=��E���K`k��L]��$�?L�� D���� P�� �o�fuM�n��qմ�Y��qd��&/�R���哽~s��럝�_�u���lؤ8�c�u-��� �T�@`k�>��A3[�t��%3��P߿{{�hC     8!)��&�#a�Pb4��!.�
ETe�,�p�n�g	�3G�{�ʢg$Pn���J,Iu�U�����Ꚙ�PV\�'Fx V�,%fk�?����O带z>6���:U��-I�Z�sR*��05���a ���=��t��%����|������     8!K�J��T�"���L�	��+9��V�1�~���f����U�߸����cU��|��J0�n4}��K��6�!�>!�;����
���^;�XǊ��NC�9�CS�~4���"9�S�u��
��x�J�ՏL�}���.��P��=��Îw�<e	�����"D;B�ԇ0@�P�e}`Xoq�w���I��*�"T��0    p!y�Ҫ�d��,@&	�H�P�@�y��(��[��]�U"6�t�Ac����}���2q֟b *y��'�ffg�Q���X����H��O7�W �� �ޟEN�u�Y�tg=��n��b��

�s���J� �=����l�z|��{\���Fo*sT�O>�q `    !��.��� �@)0Bc ��f� JhOd�GZ��u�ƃ+�+%�v�L���=���1���O	��