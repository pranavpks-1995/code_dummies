΅@I��"p(�!� o��ʒ\'4���ba��?z�D�[�o%fM�Bߩ�Hv�}zB��tJ�
  !���E��`$�Z �C
Y�	���F��x�t>u#�{|���V7�V��T�=���y���	��
��Î�w�3�s��*A;�?�	y�맒4F1�J�QbpI %�G@u�;���~�����0�w,��Oẅo���`f k�T�2��  �!��<�4 �V`  �-	�U���"�]��=l �R�dS�7���(s����7�� �;*�(�p��4�
�����6�9/��r *���e*i@��� X������ܫ���ͽ�^�t��`K�zۙ�r�!^�H����Є�9�
�jWf����
d�� X !��H��"J�6Dk&_,@. ��$-�RIK1;�&��V}�&�LP�����ǭ���J_�[�|���ʴ\>驫7��I!�_+��׽uQ��&�����N�9�.u���.w�2x� �����U�A�`S( ����_
�!�=�f ���T�J�@` �!��P\d(aQ�Ѐ jI��I� D������eu�id�@�D�wfD.�l�J���s*ˆ-����S�6��L�rc�Wo�`k�����քe:k���4bR@@p��
r�[=�Z���-�H��k'�KH�hV��I�.٤*� �h�A�h�!��=j!���f�A  e3�6��i(J��ݶ˦S6�����J�nU\����`Ȅf:*���X�hRW��.��_Y{u�����k�1���_���,܃�=�^���q �h��@� 4�����j� d���j܌��Z����R�w-,ѡzB��@��(0  �M$��   հ��W�C��,���3H��U�l�Ϙ���8@2͘{�J]����<�Y�۟�œ:��Ԉ���j���ތ�����K܉	�,�..�S������҄�Q_b��r/��ad,�Ek��I��@b&o��8�ȟ&�@0yi�f���{\j��`-�9�/���uo����ʷ��VѴ>pi���'ӼL�O¶ U��޽D�U��g��f������-u���g��(m�i~�M�J%�妨�m�.2�K�ո�*����LYS�F����oڃ�C^�Ĥl�u�Yr�ū������y�3�i ��{B��O���z���GT���wS"l�tY4��8�p&��ey��f��}�]3���Q�G���
��7=�A�7�����J��x;iUy)��aL
�ʖ]R`�O�g34�t��C��(y��y 	P�r�Պ���9�]�����T�cM+C8!`D��GA٦T�yro��ʓ����o�4���񪖈�)�Q���@�Fj�;~[���l޷�f�q"�I.���2K�*��tc�b����Jx���(x��u�v�vڭf�ʋ�b�!�\K�	��
7w8�%>�&'�H��$����{|4��V�?:xF�����L��g�R��M��u�T>1����c;�k�*��~��y�(|�s���s6J�z�-��/���tc��16�t�oJ�ؾ�R)�$�K'��4 8I�AD��G��M�T&���ܨ�j��QKV1F�1L�ԞE$׫�Ǵ�n��x�=�ۧ��ҥ�U��J�u���&�����B3���T�U��/�K9����Ú���ES7�4t�.��ի��I��ɒ��*jD:GyNE��ҩ� ��̦�H�M�B�E��1'	�e�k.ju�?�rW���C,Yʕ�r�#��=J�4��!R5k�=�l	�yb�}�_��R����E�I9������'����3 �k5�&�ڿU��+.���d����/�{Ȏ.���b�gt��ڴ��qQ�_r�!NP4���=%��DB��d�Y,~�{p5���(�کn
h��+	<O��bw�e��A~����Wq��E�qA�}�j��H���ya���)��1�ţ*�C:>�fc��G#!���y���l��ٞ������G��B���n�V�D��#A4ҕ�<�� \��Pt�B�i�b:>1Ü���1`�X��H7�q �c72�+�;ơ�8�[A&\�{R8���J�y3M��DĀ|%������K*�n��v�:��':��_�0{k����*rp���mV=*��p�I�,��i�6#�zy�CT������.�I�-�N��
�JD3��ֿ�ܫt��w\3�;'6	�!�I��:]x.Ր����\���\��mv�	0��z�3�1J���ڿ.~�93!��T�o����'9��:�{�U��u_W��^�h/}��xb���i�{b�^N���x|G"]gގ�ෙIO����{R�=k��Z��l�uG��B�cf��
���,��Y��>�12���S�	���׭�dOwq��p�-x��u���ޘ�>GDi�L)�ĝ\���Qu�o��PM��t"�Q�N��e���FӖz��EI�fM�=m��C�ӦS�?�1�(WY����&�^}Ǡ ����w�e��J�Y�����Q�DPI���s�k���-�HP4�SI���	3�?u������tYb��﷚@6���5�g2��K&��	��t�X[��e骰��#K��9����e&�+�+q#�+�5�ݣ�_+n��⿯(Q[l�g9D�α����`N"����{-��S���Ŝ� ����a�d�M��������%�Bo?�����/��@�j]X9�\P�H�(E�ΌU��-ľȥ�E�opE�O9��1ײ�D)hv�5P��$���@�q��3��q��?�<��=��v��N�^i�q�)@�2���
g�����&ٴmڮ �uA��l���HM3l���DOcJEz�?e�RP����7=&���[����EI���/��Vc#ʛ ��\�夣���U�7��2��pT}��y&Jˎ;n�LF�5UN"Vw��*������`Nې�R��K�5���9Bbʻ-�䭳�;Fg e���;�=��Aa�q���ܺ�/�z��t?��om]��-C��k�v�Ǜb�X	z_(ʝ�}�At���:|�����}��G�0�����{��O�(�e���sd	k�遗�H{
���mG�/�c����Er�k�2�x��sΧ~�@����G�v� �"b��2�Ɋڀ~1�o�Z�����@�/r����A[A�6��a`��]����\���>�RM�N%�Mutl������l�# �]�����xe3�sڂG׻�htC��gh�5������Ӓ\՛�\ՠϵ���UC{yB�f� �ځ�җ�O5-.ʳ<c�;����(��x�_��Q���8��L���[k����i���)�ر[����V<��8���;'i����*�ەI����Ԗ3��$��-9yǈ���[�i�	�ڃߘC"
H@��UW����J�ּn��LR;s�.*���1�*X �RyJ�@B��^䩍%���^��LY\g"VN�>g��!xD��������U)�
�刚�n!�-"�ʃ}_����\F�D�Էܠ�Y�J���^+�a��8���q.�l�P:%t�LI�h�S 87���R��<hUX������L�۫Z��|n��+��q��ʰ����XŒ��
��_��S�,j
�  ொnO��a�9�F�/�`����e� ������=%�ѯ��@���>�)p�J������O��LKEB��rU�zU����߀�!���~��3��4��2��&�X62�d���߾�#D�#�'�� u^�Tu0��2J�i�����l��-���* ��Fa}��R�����l������V�Tb"��GU�LQ��,�K'f6'w�,Q4�C��\�0���l�
|ԣ��k�Q�$	�JUy�"�CZ�����d	&�BD]n��A���  ݉lb���iZ�������|���E8��H�v�.<��y�8E�k�}s?d�� e���01@X|͙�k*�ʣ�R)���^~�^bs�v���H�İ=UqN��C��x��Ԛn�qokaTN�֝*M��X���(s�����
��O� O��9�H�S>�P���