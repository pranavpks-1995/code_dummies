g�u��gLӛ	�`���!������
[�&���]��E�����wJeP��Oи�3���'E� ox	gř�L����g�L��"���Ҝ��Իpg�:���	��E;%1�e_���41������9&		�.��gg��W��`u�UG�\x�4'x1]V�jO�k�'�M&­�eu�A�P&���Hr-.��*ƝX!Y�3�����U�e7��{v�X�ȧ�*�Bf�!p5_q�G��Ł�^8���l�<�KW�6��R�<<s�7��킒�3 z%o�@�(7��s�(�B|$/-���E����]ўwY(�s�>W���\%�0OI�_P�6�gu�h�u|�C��r�A錍��<Sc�&�ۊA��;�S�Q*�G��I�0��3��{>��n"'o0��a�1�?�R�84��
��8�
���B�O� >��;ڃ����̏h����3򌧳R�$$2A�,�hT�ـb�4�ed@���h?,�Q�qK��=?^@�$|.���v��
�D�(�	g#�}�n˩ Y�+q�w��-�o�̾K��K!O��j�AN�R=7W��S�m�ݩ�,��+�ahG����  x�H��d�`�d���ԑ�
���<�ޔo\݊�k�)��t`&	�� ��~�r����������VJ����*Gy�"��Q�龧5������<K� ��v+��4� kI���Hj�/<i�'����]JD��k�*LWV\�+���)��z�qtU7vUW)ļ���Iܡ��@Y���D@H{�ѲG���]�2�.�D=X$���{���C��E�G�<��R�.چT� �%�f+�NYr˝�iX�"��;�llF@sqᰭ��6��&0�묟I�՝���o$Z��6)��r�H#�g:���ۅ"Q��6¦��f���J[�55�?�Du1���2���VFqݏ�ocm�2?�Q/Uf�?���Q��i
G��f�׊b��_n��c��FJA�9Ճ�<oo�ȅP 0�뉬L6J�Nܬ:�Zzn�,S�u���� �*<��P�Q7@�1�z��hQ.�B5Jk�8�:eq�L�9�.�dG�dF;���W@���&pF�0�[�Q������@UuG��z�~0�I�Kp�GV���ޏJ���#/���~�mm��ĝMԬ�����%;�1/[��:���	8ܕc�bqD����h�=o#\�y^$%����LT�AZ�,���9L�1��+�c���+R����Ӂ�u7٫*�JJzlT���hOSƹ��[������>���s�ɥpA��[���쌽 D��^\)/��U��,T�X�i	U��w��w�{�-/�X)��5��`��4�x��M�4p��ԑS�1�P%����9��+zQطh蹴e���{�
5fz�kYX�m��QT9���1b��m8�{k�q��VD�&��$��z� �;:T��jP�3����*�L�˒I�F���˓]�}Z�|�a�`�p��5��*֣Dr�H  j�B%R��c�qέ������"���'牠�K[��E�"�`��]�/�7���s�m���n�ew,�{������(��OC�1�s�U��q��3��P��]���p����ӳ���6���!�<�-Λ�v�g��K�a�A�N�ю�a�����
�����Qkkz��%|r�G���0_Y\fi�;����I'U��R�v��g�����}�X�lm���=����^�1�e��Qupٜ�m�Q�`��4ZN��蘖 ,;_��>#ل���R|���g����N�|�(l)�<��|S�>d򶗙J 2A����Q��x��V�Ʉ�||����Ʋ���dbe�2E���\'�w��H�Ę��� 	�b⇼���bNq�?�ptL�^^P��1h�i�$���sc��
��j�&��k���#�J���a�A���`�L�
�,B[�':C�PM��5YV���_�_ ۽�0f��O��8\��Sp�zʠ����"U��nA}۫��f����q|;.����������N���y
��7��?Co��8��%E	�i%�*��I��E�}(����#��3@]q���P |d�N
��]�N���2���*�Cnh.5U���҂З<1�.����bkhHA�n7��J|c�c�!OMS��3�#!V�n��@�P z�j!��/�k/u���W��Mٗū�q�K	�y�VĂ�0V���TA��a�Ϩ]����K�!g#��(| v�*l��J@;$���ycd6L��v D-�I"�j(�!���@���1"{:���,H~����"^���v/�B���e*���ʖt
	G�_�/�I��g�J꾿���<�:����:eJ���J<�Y�O��v�������JQ�z���B�6 �tu��X�4>���Z~%y��'���~��'��>.�>��B�7�~�~��Y����\`͘�+�
�F��`o5J�Va�.�M���P%ȍˢ�uܺ�9�7��@H�;^�>��[8������ۖp!�k��G�v&(9F���R@F��\L�)C�ef�g'����t���w�jT��Zd�{��q��屎L?P�U<�P���{rD_�Q+5� �r)L���ǈO����ITأAʁ  � �&���,ta�2��Q���I�qE
!#O����U��8$�G�H��b�xH�9)l��,��ЍJ���X�9M�\�҈���{������:FNT�����z�`��R�}�q��s-�[�&�{sm2#���%���Ur��X�x�����|�bh����J���d�yN�'�\5����7ÀC�BzR�Y7��$�~�vv���٪"�Gl�fD~��OA+HeZ��4@��Ju��ϡ-J'�Rū�� �����*��.)�8�yde�J�]���@��\�C,���7��^ĸ��0�LcB�˫�!*.p�玝Z��~�K5��C��f�C�BۜR'�����y���΃��(e;,��Sv��RV�@JD$�b������zbD���o'��WQ�;>To�����|���Tl:�a$%�#�kC�L����2�A؁q   � �b-W����J�9R#D�r�s$2#��V?��q PBW��9��<:lXo!%�~�(H��";\��U�C�]Yl�=+�-���,^s<_r ��D����O�-�4C�u[V�������F��A$��n~�b�b�	I�:9�S��T��O��-�^����U^���2-���󸲆���o:�>��zks=rH�����vF�{%�MKՒ�?b'���7 �n�뼻*�2>g���-�g��.���t57u����9q�;�����4��%�EbZR��S{f���X�d�{gE�l��3W^����g�Й׷{�Y�Y[���ИŁ�+��0�U\�:�X!|6��b-�Z�cH�W\Da�N�HA㪩*�0�y��a�9�G��~�l�p(LLc�|�-���@��2�X�ʍK��i��_�l��ͨ�e�8լ[�����7��,@��	�yӒ�e��� �E�:��������!y���	& H�P&��`���~���+v��G�D��/����ws�dg0���	�Ei�����PL[`!9�0�s@��5�rBZ%�������dn��Ցm��3�D�\��܆���V��t� ����-�-߇P  8!���A	Т0Un��Z,����  A)���P���؊����/W�p]��pB���Vl�]1�F�u�:�.���t�.=%���HZe`����oq�e��]����&��S�3����>]j��wEp�5 ���  N��٤.�M�'�@  �!�*��C���T�,IfCz�zR&*�>�����xc�m:�ׅOkp �P��:n;�<zNL�dnSV_�|&��Ay����5���Q��-�_��6�v뚬�}�kU0(��l�Tv_º*��8Sb*fu<&I��x5�zA�L�0�Z����PC�	o��⪑�u�Nn��H�  � �!����!� �uU`Y��<�LL2\����%� 5������h����Q|H&0��O��<&yH*;'��Fx`Z�k����!�=?�kY)��(R��� ���|�tW�f"�� ��@xJa}�z=a|jA��U��f����v�}����H���P !��.�� F�6���]��C��kVғNJ��8�f�\1�A����v�YĴP�}�xmu��.�g�+�îԾ쟿#��0aWzPrD��X�O0W�'�-D �@4�ѱ�'��Km��}���}��n¼vr:=n;q����/K]��  �!�a�&*P*2�p_-p �Ml�Ĭf���Q������Y�ֶr1V�8B+Β�h�_�m�����/,���Ȩ�p�K^kG�
L�Dy��^�Unn��VįI��	g����V���-3�@���m� 4�*��Z%Њ� �   �!��5
�# �b!!LS(u�0� &WM@c,AW&�ߪ��z��h� SE�EP��"�*N3��˷%���G8`�� � d=,��y1n��@��[i�|^oB�F9Ɯ˛���!Ie�S�k�v�V$>���{�'E!�h�n/�HASją�b  `!�
���b�b��UHp�ZH畁�x�n^S
%C*�$(½�3��F�cFޢhR�j���$��Z�1���5��2.�
5�3�`� hx���ZVRO��V�ɏsp�(��P�}��΀&�!��ZH畁�H]S1�G   �K��l   �ӈ��W�C��I�b�~�(�4��Tm�CT�+��X�����9��b��br�3q���_��yq�&�˝��9��iQE��n�����6v�ni��gA�=K	,葥�?:��N�c8@B+]̖���(�Q�����,�GF�t����[S�(y�9a?<��j������pU�'���l̅��l�J���ɓ9�J_�C,�-G�S�|��4n��]x�8�Lu����U�!E|�T���0Mmfbi���`��v+y�v=�����p䍞�o_&R�f1{j�ҫ*��"�.�)����N�T�0�y����To�d
��Z��+���a4\�P�O��['-�>��������l��V��kO2��!C�cgE�t�NlI�l��B������qH{S�^������~wz��G�yE�J[����H7��Bb.��C?/�y)"3��83?�p�t��#ҭ���mO�A����S��T�"�9D����ș�����ҁˆu����uWQ]�F������Q�N�g��� $�5@�c�������[xp����J��#Yi�����j�� @�C,ћ���+����B��b�l�v��-�+��l�io�)�Q��*%������?rJ����~U���5�14�pDQS�I@�#�4lǧ-7֩\��TP����B�`���ER"��[�#A".���VX��0�w� ����)%�栵���
����ң�A��f�V���Ev���O+E��}�#h���6��SYȣ�'��mV��`w�#cU�9���bT͓0-�P{�W%D[��3U��� My�}�X~Aofw��
&;��p�(����5���LR7:�_|  F2�1�}��JB�`�௏�<m��)���g�x�'�Z=
�L��)�zL��N~R$�}A�������|JnşϹ�V�3���JMg�{
�7����͠v�:S&���X�07r::�x*p�?��"�^Hו�ռ��0� N��h6��}_iˁ>�/��B#Dmn`s�t6~�����[U�(}"B
5>:��o�H�j��d^ ����T������GƤ3�'i�@�h-�v�Ɉ�|1�$�`O�zw����u����F 螤�l���YtK�A��%/Oo�FVR	R��1��;��n�U�ts��Tk_nf��K�u�M ��E��CWbhڠ�n�<^KW�$^	'�sd��LR3&��[-�}��m�	��+1"��A��7��\�C�������1L����-�H!}�F��ť��E��l��;�MA�N�lwZ�z���� �̀06�"4S�&F�_�:L�0�b��̦�?�{��7�0���J��X�Ґe	��k�n��h��[[x��"�:D&�:��*JU���b>62��
�c/Z�>�B�~�n^�r�2���dGV=�D�?h���