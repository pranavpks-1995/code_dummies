package probaData;
	
endpackage