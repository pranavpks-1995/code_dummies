\'n�A&��#�N{6a�(�3E+t�&�������z� �Y���Þl�Ce�x8D��^̭j�*P	�֍��,��,.L��n�;0��%�7r�#uy�J�O����������SH}��M�Ц����J���X(�;�j=����\D�rx{,��N�E^ˎ��'���l��7��#���͜�	t��u�����I��$XP���'kۭ|��qb-9��6�dX�OZ��(K�JX�wh%N��?s#�{��9{�:�4t��9��=�QvS�k�r$Ȏ>mEAj7߂O���f��H�d g7җ��7J�7���sxDϑ>^�^h���W���@��j@ı/��o�e@���:�z�Dw��t0Ԭ8bquP�A$���?ה�u� ����:84b����`�-D�ܜԿP��K=f��3�|8�\b��ߘ�s0<� <J��G[^a��N6؎Od6q��
-
�"I��A��۾'2�8F�?3Ii%��\��蹿ܪ"��Q�&����Q��5��s/1�/�Fx�4�$�{ d��i�sȨf���T�pDJ��h�)*aHt`h��sӛR�D��)��c��f�òA*x�DDY�i�7�y���Ul����#/`�"��2����U�CuAg���X�6���9���&Zf�q�+%������'�s�1�7����	�2L�E�c�0
n8��4�+�{�|ڑ�9�]�	Mc��<��Q2�����8�mӈ�/8�U�@�$l�Mq��4�"K�߈��v��2gF]�Ai琐�e�0�+�~��u���$=��ː�Yo�#�Gxz��6�ߞɡyϲ,2"�:�E7hm\��H�3lT(ƠI@9�;�n㚾g��5#"���[v�ˤ����^G��L���UA6����gH#C.W�Bj|�1�gd7/��(;�҉�l���c'����|�)�%ߥ��R#�������u?IN̄`�h6�	���)���2h���}���5A�,��x%,.G��o�a�R��j�-������o��+{�I�4���k�!����1!���A���  ��"'R��c�@������@�0n�ϹfU��'VoH�p��&�����*�p�3���,/�7U��ߓp�0� FZ}��~�9B�W|����R6�v�;��K��:w���
 �DmU�*!���ԍt^3gt B+�,0rt	u�B�f+���r	n��Q���j����o���f���J8E���)01@��`�p1̖��Kȷ�X�$���{�܈�j�NUh�$�Am閈?����0ٙ|5���,K2�� Qx���	�y�Xo�}tF��=��,&���e��&�ie�!x"���r^��q����C��/᪊[T#����d��q����� ��5���5ŃW�iG+�;`���3+� �f=B��M%"ט��q�,�@��>'�������Ѿ
�!�6�m�����'�X�b6�A@�>  8 ���U�y�IL@H��D��ޔ��=U?q[RJ��B�(�֣��YYSF�<0w�ỬB��:�TB�+G[���#�>�8�O�b���P�و��i�����Ԝ;I�s�R3��6)���*���[�r{m݁�G�}t��8�ⱅ0�>��DI�,��vA�v��Kͩg�d2\B�;yHG�+�d	�2�D_p8�+M��h ��uU�u�cp��(�aUf~����l-q��h+@������3�3h�@ivG� �X��B(�X���C����a̿;p��!��Zd�G;�n  }i܊I#�՘�AW�h   O ��u�y�JTtpR�����ѧ���zW�/{�̂�O�҂�J2�8<//��۴F�L�[nn��S^�����u1����!�&lc+7~�±�3�w�x�NT�ONUW���p(_��uΒ�U([�Pά���c����}��pl�POxؒ��C�X�SŃ+�J`�l@�Ֆ\�V��M�;�J�\�@l%B}@#�G�J@�q�'��K�{���֑��TN�7�Ѭ�PY��������4��~���c�O=��A �=-5��f���4ЀXZ��a/�w��T�nZ�:�^O�\��kǏgqVøq�.��*0Ӄ:S���	v�� �{�N���@���    � �B-����sJƤA$@����= �zʋcR��{,܃��^"�e��%��u
Mlږbw��P�?���h�N��0P��p8��>�-rw��j�