d/q��!�蝅�\>�>^���A	
��R�t�ǋS1��>���NͳLRvz?��^:W�SAE=�.n��9��n�(6�&�\���Ŭ��
0hX4F|t�Ě�T�3>p4����",�J��hr`E>/oT2�S0�v�?w�o]��o��ޤ>������d���J�0�x���K�n�%d�ߵ�\ܺ�J���r���ꮁ�5��:�.�f��YL�ݶgU:S�I|G��8�7����F����}��H�O�2���j��-�����Бs<�5a뿜:C4�>��p�(ٴg�΃5�hW�D��K��V��@���.kxI�z'5@�!��C^�E�;6ޛ��I�6����#�8�Rj6G$ҋOeՒ�V�y/�Te÷���
Y�b�%)��12��L즇�{	���� ]T^D�,(X�~�[�����7�V�3k�N�0��+S���5�[9U�T,��p��*���^2b�ͣG M��N�J�� �=�$�#�c����*���j��3!�����V̂��q����9ύ�ڲ���ko����R,J�h��gd�2�FK�[>H��䶬~b �R-�J@k�OS$e�rǀA�2u�T7zBaKKw��wR�.f�v�����s����I�q�\4�.���ƅ8f��N�3
Lĕ���i��!)_���Y�a��h#��g�Ė�e�~��^����"��&14Mg��7����M)I�Q&P�'�}���8XφhY�(	�m��Ѷ��M��ޏ��ˡ������?���}�1�[�O�uҺ��%y�h���Gvy�^��g����(^�����$�{�?�x8?��3��%kЕJ�;,���=��ͦ�n=�=���[fI�>���<��:"&�ݼ�)��\�:W��*�u�AZ������=��C�d.����z
�is�ôMNr�9��\ܠM3p]TИ���Qx0t�LK���?֒�_�HT���&Ҝ�UP�bfPio���);�p��)~I��x,�|�6��nON�wʳ�Hz�7VN���g�Ю?	�b�J�d,�0AD��+���Is8����֒2�r��fL�7뽯��T-?�*A0ݵ�Y�i0� �����d�ء �s�ˀrx��ι��ű��}a��)��U3[|�1#=�[?�Z����i���]������q犣C1�ʸ�^d�.�� ���;C0���w(m�J��6ʸh��+��=�9�1b��V��Yq^�:���p��r<����ݹo��ڢI-�j��<�G��������%�eW��y�F����#H"s}�N��y���(����M��>�V��V��Y�ȍ02�{Ѱ%�}�