0΄Ct�Y��t�-V��I��䟬�~G�ᑋv�aP�!�-��d�=��Wx�c7���^G�q�'
/� C�Ī�|�����S9�i�W�*AL��'�hq!�u��V`�,5)�x�;�˅ڊ4��K2���x��G3ϝ쯻��D� <��'�A���
�wW��*v;4��c�1Q+J��J,���؎t�6��A[R�g"~ЗUE �c�_6,VaL�|V:��XH�&����Dt�go#��I7�R�7+�H����X�8�f�@)�l�!jn��a�������ږN�d��>6r����Mn�`x$'��4�s<봮������j5��=���k��\��7��A+\~����xX��s�|�@�v0����X������uH�:��8�Ȣ��s|�������a�ry8`������X�S��ަH��*��<1`և9�R:��%w��.v���,7�wԛ�'���
�V,��WNe{��M�>��p�\W=�� �H@h:X�jM�Z���#ӎ'B������Q�V��P 'C��`v�Df#�L�@%U�c�j,GԿ�s����
o���	���ՅmF,A�4^�����Ϝc�b�%�k�4���B�y+4�5�Ᏽů��RifKfe�>��OA���*������7����{�l�d���*����'�7�}�ЛϠ���4?��jsIu�����|�FX�;�G��uE��_�ɣ���V���p�t��y�`������:�BW�J[~v29���z\�LaD�zj87,�}�K�`�-���<������OXsl6�|>7c.&.V�⃯�||stO�9������T�>\�V��y׭��]݂�ݧ8x�w0���G�I3K!�cP��t�Z7�:�Y ��e0 H!�(i����К�G��*�=r#��y!���i�I���n�Z-���&+��_UxFԱq#)a�Cj�r�Sg���9�ʲ;(/+C�/����
P>�P{���z�� ����h���Qu4QF��=��o��q�3�Wg&]��>���C��(9�;�}�R-�i�$�㯙G�2k�����kq0ב*�z-��K��@Z/�0�-:#���9����qf,�V����'[��H`�Η������11w���D����o�e+%$�-X�}�21l�t�|�	���TDpU����Qz��7�:V-��|X|@4�$wW
ZN��IK�L�x;|	���������}�.�Ul�N�V��86.kҁx {���-!m]��E�o���$�/�ӛ�ElJ��弴���R��V7�}a���]��%����ѽ���ظd�H�z(7(���P\���o��s���C/ƚ��޲���	�A�,��r��}I�n�m�աD3���y3�����C��3�6��Э����<9ȭ���\���t�C��P��TF>�Sͼ���RI��_�2���W|�0u0nh�����o��8�#�19��g٠��u:��l��E�8yGe3��غ��X�9v6Ϩ�/K��J�T?/l���0>�p���Q[���*!
TP��ZdPҧ���b��n.�x���MAq�_ۂgC^�L5hy�n��!�=�d�Ա��H�B�A(���ͷhp/m�~��Aʗ�d��V�*��K[�NnR!rV�E#��  �'R��c�I0���A�5���@���'���s#�3%Β �/1���i~I��8���qs�t�����3�y�	�}��0F�`���Ǚ���OU>�)h��v�_��~֊1���vg�j̍�M0���(%�վ�,2�Z5�찜{���=��X��5F����f�љ��Uؾi���k�V�.l�.d���S���k� r��i�ؖ&(m�^���.¦(��Z���w�����W������<Bu�#�=ѾA;롺a@h7	��F�MA! Z ���
͋?P��[����AR���,p�#�λ*��9�d3�|�d��]̗�
���[�}�sj��>^���RV�ùɒ�2�	����$ f�3��8��1� ��ᧉ�������9��aRZ�c��8�P�Ե�p!�Jؿl.?�.c�v�m�c�CHm$Ԭ�~"����7��F8t��4�k�:�肑�lۜ:���{iw��$3i����lЁB�@�M����b��A�v�iPN�*N���K�B�oǉ7�� ��.8�����s�8H��>^���'��W�;�l؅�dZ\Ȏ�K�������Gl�F��N���~�Ә�N�i�Ns�V���9W@�1�UC��G��MLw�~O�#p�b̎߀7�ԋ�Em��u*5a���?V]��57I*f��3���X~A�^��Ӯ�����(!�r����?��ߧ/O/�=� 06��e5)�<�x�Ų^�72�?�O�:@k���'2�m��5(��[ϳc?����ac8���<̇��� ��\{c-���B�-o�̡�M/����ЏԂ�K�y�</8v�50B��򱸍MW�h�GG̲�z��U�ݿ������n���(Z�c��Fo��;?�E��e�e�'> A�5;mZ��s8m�X\
:��`@���6w?e`@h�����5S��?�J��T]S㾪&<��ch�!��L��P1J�Cy8x�$KO�퀃kf�)�DP�z���ܚ�QZ�	)�ͤm'�{����-a?�&�����v�Lˇ�,yuڨ_,��@W�'�	��>�1��B6�)��K���1t��3T0YAp��dd0p��YD����.� +�dŁ|�!����B�+��e��������i*�Kq�!�� y�ӣ'����*?���Ź�AE��(%.���kcا����7��ߤg5�.E��I#�
is=O��,@@<�^~�cn��g� 2u�V���Mj��Eۜ�A�l�����6��ȫI�=�Mg����r��x`�Cz�=  r �F�U�|�6�%4+R�����X�6��P�����e��p_O7/�����2������'�v��#Q���1�	�[�l ���Fui���W9A�\�JnT*�YK�����{���`�NVW
�R���(j?�f�;?Ѽ�8�¾͏{���>KZ���۹}��_Ѥ-^d���E/���e�-w[����%�fΗ���t����/��J���1����P�"_�>�-q:�d�6조v[�=n�Pz���9�/w��V1�R�j�O[���+��m���4f9O�J�g�k���S�Sf�W��vM�y��Kp_��C��0WZ�����yMG��O�:�������C�͐}c�𥡐�2���p��Ҿt8 �0�}P�s�#^��{
P�k�����-�W9d�&��1���D��c��2C*��9�Rb���|[�|�*���Q���PHmM%
^^ܾ���0�N��ws:�����%@��3PQ��\�3��L<�����2���f�w'N>�rW�ý�>5P'ﾌb�S��]4�lBB�Yֻ�!�G�>XZ|��sɚ��ZN
jhMZz���B����s��@�yӤ��ƃ�7�,���*rm�}���]���GM��}bΫ����G?땒�y�ZR��^�BCˣ΀Ѭ��n�.�a{j<�)(k�� � Z�����z�Z��G�2-w�����Ne�Γ��,=�~x���4ʎ%�K�^�F����U�&�������4Ho���d�AL�*H�M͏AIƴʩ��Ҥ�����]��&F"/3�}��X.״?X,��umυ&]���i��O��J a[�Gv�Y8|�)cvo/���kб@�Q���eI
�(�C�f   � �f�u�{k$=E�hs����!�����Kd��A�~HKCY�F>�-5�O�O���j_�L�#|bQ��V��N��t/�b��b�D27���j���Ox���zu0%q��0U�,�~�~}��Uu;L-1v�{�� $���h�(x���K�v*H �f�E��6*WB�d�:,Z�Ɍ�|��xG��GH���<�F i��,��	��*E��h���!�1f���0�9�P
�q�6q^�i��M��/��.yЃM�]#Y�#BAKx�Z۠�gH��ʷ�xxhA�HT��k`���� �9v Asc���A)�`�@����a.�
�FG#WM.������C�o*"h��29l5@q"��xZǳ5�4�Kg�Ͱ����v)�b��/"B�E8�@{��FcQ>��{lC��-�Y3�yk�uKs  %��pۏ�6�(����ћw�J8yG�w��ntc_���%��8J-��@`	��M��zJ6ĵ��I�C��L��x�-(HY�gmT�mu����C1��.�V�bn|-�Ra�G&x~��J�C3��b�Հ�qhp43*�\��4���~+{�L�8ӓ&N]i�ZkZ)�4�ʾ-�����<�� �oכt�F�&���,�K�(۫�~��P�/��gq�@)zW�u	�+�f,ʴ�z�����N= \�&��M���ϟ�ƎWGiR-�*I<��HƜ�a�t�Eقnx9�R{��_]�W!1���ni��W?.��(%+A�?S�7���B���   � �-�����N�9���2q"���CؽifM
Ƣ?�2��m��sw�M�Z��v�B�C���>�"�s��3�A��˜�1�P��`!�3ක��UM�|�V��r�S]{�_�؏9�~�w���D�C��|�g����4f�Т&�x㡆ǻf#�|/|0«1��ݩ�O�@�h�*�_9x�(5�G
��+�S�N}�e0�I^��SD]L�S�
����9��#'ܺ���
�ԇø1zو��&�T�^S�v��Iy���Y����iS9LW�Iu�i�I�-V��r���@��	_��Չld��WZ�OX�~�S��U�ɧ�l��j���=��;�Yb��i�!  n�����@Q�@4��h�G��O���)iS�?`�I�P�G�]���A�q�7//�bJ�I��海M�E��	�.]czO�����֎4�2��ʿ6��U6j�Ǡm'�]��9R���y�a��U&�q��4�"�!g����0w�L�`�Z�7�$�D�Nԋٿ���1� :&?����D�L	�B~�w�Xᯂ�����
����v!	;7Vo.�yDs�OtӴ�ޯ�c�J�omj����~?>��4\2�D���5���>�q룳�w�?5��j�z����E �d��������!�����7V ��p@�X�}(C��U�"!3o��*�f�i�������$	�5�E54w��@y�:�׃64�S��劒�	������=��i�9B܈��U"��	�0�(! +�v`�|�%�E)��U>�;�<ҮP�#��U !��A"#�PWyBL�G@"� $|g�J�dB`�X���B���K5�UZ�u�:;lڵ[kJ�XpMa����T��9ݚpWBKE3^��\��>H宠`H �S��@� �������=[�t�;۵��Z��bѡ�8!�E D�<+dCWlgV��mˆD��W�)��o��C&���
�S�S�@u�ދ\���Ͷ�/�a�#���;5�].B�:>z,�\�!�{ �t�o�<u�n����U��W#7�(��(U��By��� �o���=>�+��+\zj�4��ۤ*��Q�Ÿ��d�!���"`�DJ��PbX ,�f�D��s���e�Z�A���q�&�M-%k&ū���B����,�@Z������RS�t��c���MA�Od�jF��/�d �-a�Vm���wI �0	� |e�}�ô���]T��r^�r(�ڹ�@     0 8!����%"�%69`�`�V�t1<%�;�e��\�u��c������w2_~�/�����$�@>L�~�^o�9�;������/�Q%�
��� [U�#dB�����A�(;̣���yܮ9;Љ�aѠ��5�|(�y)�ޭ�6��u�,�� `     !�I�!L�ѽҕ,C`-m`� �A .mK�F�����T�v�Y=�G���u9�s�o�����U
����a�f �߼Ӻ9m�n�f�(�Ku�b�m�}\;�y�����%t���> 5�,�y���t�m����������N���� �    8!����E�A����@xwu�f�Ŋ�DrڨI�*�|+�nճLw�'/��#V��Yͨr�S[`@�7���Ӯ���CJ8jC�$c���P�¬��N��˗��RR�2�@A�0 xIC����&uND�o�T㿼��ǹ�  ��!��5�&�U��ʑR
I�F� ��Ԡ�i5���
b�fJXh�-7�Y�M����RE՝�Lb�� �x\��4�/��;�����υ�\z����\�Q^�<1 }�d�pHaUR�<�@� �!*� ����GG_���Z/����0��b����Tp�T�     ��Q��   wӘ����C���%m�����k�H����ņ���@�z�G���8ѧpxB��[�g��N�\G�GҚ=�Ag.���v���h�S�}]�_B��b`��e����8N�/��
���N8�=� �0~{��v�I���͘�|�([����*���d8��_*�Xb�k��A.q0r����Ke�z,�w�8����eo���F�X1�2���/O�#�1��\���MN��qB����Q���lڑ]'m�B�g�7��v�ob �p��"�^��?zm�k��a���j�J�V�Œ�,N��D����<��������`�Cy�)�P���G��i�®�,ͅim*��Ǆ&�V[%7� R��� �X=�5��N��!�-��z�wl@�NPDs����niQ���܅�/�r�:�Ig��gx�4.�#I� B�)1�^=�K��P�b���5�T'����`)7׸x]��1�N����td ��a�}��F$ak�2g�B�@���D��#����V�s�3�2B	�(|uK�`�!�D����7nQ$[C�1}D�l+
���i(����V���kO����I�����y|�:VL���K�R^�?���-���se� z�� ��9���r����hB2^�oIg�jj �:���L�7i���o�����&!����|_q½�g�|f�Ĩ�M�>�]fI��=S�f1��Ӄn��0�ߌ���[��[�5��$$|��U��[gTv���D���B\�F;]�����Ey\��>�����<.�d�O�F��@���@����0<5'�|���4��4u/��c;.g�����[MǙ�[?�oB�A:>�,y��N�Ã����w�Fⓑ���ҡIn�Mp�Z�RFX��@���pVW�R�]b�w~�ԙ��PX|���/T�J���g��y�r ^W1Z����] p�݇�l{t�����5�~-��o�_ ���y���ͮ�#��L%�Bg���u�
d�(�5b$�ۄ�
��`����tL�:���NF�ϐ<�=�����'e�J�k��ݷ�c�9"��E'���|fT�
y��H�ƒ5�N��}�H��dQ �:�>P�Ns_:d��v�~[���[f�.��ꌱ�7G�`�@����X����=)T$U���vbd'����ȧYEDpT��U�Ǳn���c�Ye;I}��2%a�c�����S�z4Tt�5��Ǎ>_>�ٷ��_�cZbϷns����� �,�H2���@����'�
�`%v�ڃ��p�j��Tپg����JC���{ �uEU����V'���#�.���I�qؤ�|�Yr�z��W`�h�<�o��|+�j�6<o����C�O��K�*;b�P�B�G��/�:���U��R�>_)F��A��V�&�b��f�ݠF� �1�鴟�C�� [«������OK\l!�1��.��}�����^޹n�E�y����Z��*�3%_0�I��g�����W��-:�vRQG�,�0�ǿ1d��a�����SE��0�z�*!��n��:D�<e�$&�Ӫ��ԯ��
�g0�;���ui[M@R�q��V�t�l�q�^iH�d�s;D�7��!���9M">�_#qN�$ra
u:�Xi�T�f���C�@:l)o|�]@�B>@B�� ,�7�l��.U4As�*%�$�\iG�j"Bug�T��`.(~�]�
�&�!�=K:	,�y��)�LU�NUi�ZB�O#JT�P�����[��&H�1����y<��ݛlɿec\����GDǻ��ؽ�������q�g5C�\���/xǵF��N%%�S�E}TW5���r�8��J~�%ư��/���r�KxQ�e�b���=�8C��B�KN@S1����|@���tZ�2e��Q `0��]��M}H-�S�a��s噭2�� Qðl;�t��-��;���4��W@�K�Ɓ��v$�v�y�A��c�R̋��ѩㅎ9����[�\�UQKmś������]`��	Ģ�0q'��wd���a Y1�		��;v+��h*F�w#��q�K��Q���9`n3�����[b��j/ ~�@`��-���2`>RZR�1�u�g�@�f�a��ن�7��2��ݷ>;Z�N����f����r3���1��+��Wv���83a�I��G�j�"e�`�~���7�+u/.2��|8?�
Y�oM8�($�`�������_e��"f	J��z8e2�!*0Q���1�'P?5�u��'c �.��[u"�y!Mt��9�v��WUB�)�.���P�u�ؚ�N�yec����G�}��f���F��Y/��KT����_m�&�;پ����b)��ȇ9�����lp�Ԭn���~ka���1��� fkN*e<:«�_��'#t�ǜa��!�8�t��cӄ'�%߿�Fǚ�U3��3�g]}�?���ر*������݊�s��'�{Joj���n֋wIM�b�ϔ%���avR�����(gn�n%2���z��w�E;��}ת�h��H��v�RBB|o� [J���I��#��Hc=��Ǻ��N��^r��7���B.3]}[,�3�r�g����:���E<[ou��~�D5�:�T��Y�&�6l��$��Wc�k g�>	�B���mr��K���(ݎ�.�Dd����W��P$%B�N�X9&T��S ��޽����+c�Ya�5EL���kiL�/��J�މ���7�����-6'�������U��@�s���'����v�'gr�����e�8���U[}�D�8
d*øJ�,�^Y�=C1'��E� %�Wdj(�tJv���(���v2��(������}w7q���auۓ1V<:Y:�/L{4@�_����|1l�k.k��3��s�nCHy�
y�ȥ��&��/�U˵�l>h�SFbW�� eFl�Qsq���0z�5��s�%����Zy��vjj����R���v#�E7�mV�09rd"�ۡ�'D�mK:���q����� ��^^A���-%h���1���{�p1<tu�y���I���1���"�L�ju��9@������A�L�ND9�ۉ���4�Ǖ����mb��z m�S��L)��������1��q�6BC��M��9H�.�ug�""ֽ�S�C𞙬֫�<�*�1_1y�2�TNYs�lzvbp[&o4�Ȭw��u�S�T��_
ƕ־Pw��O����)��2���8|U�<'�O`�s>�&�ND���e��m�����T�[�D�7��Լ}�0ٌ�<6~�m��]���I��˪~m��p}p�2�����%����aA��E�.)��P������h{A�~��8b�l&}��)��+]���w�T�`d"N� sF����!�Q7�T�Q�r��������FBƽ�O�5㞒�F����)*X O��Ӱ���c�^"��0���z��Fzq�4]�d��C]U6��~ηG��h	����r�:�=H�;t�-hK��С~e�-$�l�z4�Q1)��K�Q�DB'������Ǩ�C�G�I�z˩h丨�䰖��b�>�p����j��`W�ԺX�S
��=%�=Jk��"�9�'�����Q&�����%������Ԁs�J:12P���p�ru,��(.�c�|��vU�0���P>[��Rقqx�5���9q}��8������$�a�%u�����(Uu�z���Ӄx(� _|�iX��@1kZ�=��2������,>{BJH �k�^�t�Br&�ߍ�٫�z�%�Q��=�-A���÷<���~i��^ߝ�ᅃ�ߢ�a�/��M�����cs��	�P��7�it��̜$$ռ솇]��:XS³`��h�����qw@E�{��,-?ԩ�@��ILy��8ێ/��QZ�xP8>������h�W��˙Q�&����?��N��D�.����M�u�m���.�ue�����+@��7�J��>�=E�s���L��͟����H$a��[-��F#+���]��;lpB���8^���8؟��,��fm�%W5"≏հX��Ck���1w�����P��V�ha�*(ĤG�W�ۢܘ���ۖ`�A��_�69*DN���krI~��Q�8��l���,�A,x<�t�"�m�aJm��<+���z�SrH��y9n-��:��#�iRտ{Z1Mjf_��/��:� ��0�����3�`�]m-8<�Ƞ�o+|d�G�S=�Ūe�&轱?�&f���f��d˴�͕[���n��}��G|~SNȢK�ܽx��x^Ye����P��=w�5�����?a�3���g{��r,�K�Ǘ�	҇,����S�or��˔�]k�?�@�FՁa  ��"'R��c�%�N��@�qhL\�֠ќ*y{+/Je ��o+��~̎�:�����C�;Y�F��\�=ۏ�<�%"�9�.���m��;h	߯�e����2p<�d�H!��P�[�!�z����3EnWS�7�x�G�TB��<��|Iv�Mr�E6����:�G�ʿL��$K�1�٬@*|Һ���7�Y�BO��A#9 B��\��!��c&�U=���e*��l�7�Y�_
Z� �l�!nq�r�ie�^�����WЀ���8깈�s,�����{1��>�3�GN0w�	���!}��E�7e�(�/�rfd)��P�L@<?t��dkd�Q���FI�XFT�^�zh*��ϻ���.���+pz4����T��d��)d�h0��+���3��lؔ�J3��4��m!-V�\,ǭڈO��_���=0Vk���LF:���'�2��K��sh@s�0��O��rm�H�;���~�ɗ��+A�4�Q�Ss���6ٓ޼��P����D�n��1{�1v��z�#,V_[�IN��,�Jgjp�=�[��q� ]���q���;l\g6�\ݿw��UZ�oA]�8�ט�h\��Zi�Ў¿c������{�H������3)�����=����{��
���<�: ���Dp�z���P�p��տ
!��EW��q��� ��tߩԕ(�U���Q6Y_���k �ÀEo��T'伷Z�
Y�T��x�5S��nV� �I����������5"�20��)�FhI�W������[2ԇ�H�nwFyN&��1N�b���w�ݖ�S�:�K�n���*��^BN�\R'���J�������MX�LA��EK_bhT��Ӥ�!YWD��}� 0#�3*lP#�}�}�JU��a� yWn��+7�`)�n[��z^kvO���D���&Ǉ�X�6k�y��*H��q��6~�c	.Z�<4�"9��8_[�'>��v���*��Mlqe,���^8�dU@)�a="w�;���ut�3b�h%a��)�"���f�FW�v)�+�� r2^~b��G���)����к�l3�5�cFe��ɒ��\��E$Og��9d���!�)y�c1�\(��ߎ�k��r�`�u�� ?������dqa����r8s�F�f��e�n�~� �r����tJi�eu;���UOaB3��u�
p`���8xM���h.���.����嵎�D��l@��Pxl��pOlF���x��ئ�vM["�:�W�(G���W?D��#u.�ۅ�3�M���K��P�p�j ��)?�P�1��4��9�Cp`8N�����h<�^��� >�|��lԴ���� e5l�%�ˁz,��a���� p��)�Y���m�!0^\eJ/f�����3d2��q%>���u�I�+N̆\��y�-Jp��J4$�s�ɀ����3�
٨ۗ�󠵌h�Od�G�An��9�,U�xAb�����w���|�F�{�)���h�֘��K�JT��D�=�~�m&`�g)�w�Ae�8��G�Ujc#�l�!�Ő��-4��rg���H육��f]|4�m������~/�C�S:����o�s����'��W�.uNG��I�ЁBiP��b����|�3ആ �ma(,ܿ���f�� �l��;:qr��A_I���`HL�,,�pԾ��]�v�3��L��R��7B� �@��y\�C��  � ���U�{Ng�+����@�JB�/n7����e�~��>��=�&��J`3�*z?XN�;��o�X�0��"(���=w����l��)����
��v�rDV��;���19ٙ��1�����)E�x˨]��P��1��צ�iZ4^�����@��&�֏`e��V�Y�A��DǛ�8<E�uX��7�}�+��U�= -���X��~&��ti9�N
�L`��c`�l��y�?��Dů������rnt��ŪE�r������Ƀޑr��ԾH��B-�u���"+��~��_l��Y�c�F��2J��?�@��zL8-��l��i.;���	�k������g�d2J/L��X���X����lq{Κ|�X�`���w�;|������S�D�������?{��^���v31%��7x�']..���`���2��f�.��^�9��/խ�0;����{���(Zǜ�A׆x���w-TK��lV��	7�57W��m+K���'��y� ��a7iW�(�����6�|_�(�9��12T,�U=���\�jVY��$F��y��u�V�KV�����K���p@����pT����@�6B�cb=�7��	j����`Xѱ�e�ˁ���P6ؔG���Or���i�E��SMW���'��i��;S���]).Ip�*N(q�:)}+9킘� ��#���C��b*�l=������"C�j�A#�T4�p?IPIxp�b�L;7��,Cz�����ѥ�.��[� O�Oj	���R֫���w�+�T'���.ե*~\��>�-�)��B�֊݀��[�'��ӔV�˔���������>ӓ����	6I�co�c�Ͳ�&�g#a�R�z	���C��&���v��N��*M-��@�D�7     ��u�xM��Gc��48��c�%�.|���ZþS�����'����>G"��l���E^�c8Qk�D5Jp5}��fF4vo^��ʼ���xoH��e���4d~��oU�h����s�'�����(�ǍZ�ч%4��/}�'+�$���jn�3s�-�Ǟ�a�����j*�B�)��z��f��!sM1%�ۺ����rֱˢS��CI�E���YR7��{`�-�>],����&�|����o�N���Pb�����08������D�����G�����+)���y�.Esn/m�0��3~�q�ª��6��ʡ+�/�J�p�X��j���Aoj̺*%W�o}�X���(�P�V*�S��`���6�Ƶ_2���#�x�#�QT�tx�P��P�"&:����/�뼏�%�{���3�C�ԑ)X����4���t�S�������	_�dp�{4>VQV�C�
�Лh4�|3r���F}pDI8�����?8�w���m�����Sm���BF���u�r��A���y�	��x���ll��V���r�=���~�����a�m��*��v��V,�6�$N-E�k��q���$���Nū�?�̏��e����,�I�č�7[--�|\�V����J�Wx�}��1��Ht�Mߦ���.�j������w9G^#�LE�'��0��kn�a��M�Df;�F��R���Ve0�?�r� �A�w�/�JNVV��F�Dt�?�щ��u�,ְ�+����*�R���\���e࿣���٘c�����Y*�ΰ���p(Z���\�}��?	D؏��e0�_�o?a��+'�)]O��RvQ� 0����܉oǠ\��4t�|W���	0�D�1u|�iz�rF��Pͺ�Nb��uᥖ�d+$�μ�ഩ����2?Q�K��Q>��וdl�U&�= m:7cJl�M�$��e�K�G�*��
U��u�E:�7���p���
n%������s�C���   � �B-��������*-��)P�t��G�Z=�q��yI���%��x��>�f�@}lC�ʰ`�NF7�.�1�ۛ/���|����W�����940U����fk	��,eJ��|l.���,��]�a�}ic���jȕ&���Ӟ�4<W̑	YJP�}�ˀ��B�l��y��}Ȅۋ�k��G0�P�_\�U�
�{b����/���A���kb��]J��w�}~��Z28� ��mp@��I��9���PO��S�쀓A�7:�����C���0��\�qB<�S�A2:*H\Ѕ��t����˚�O��7���7U�d�B�p�	 %U�{�1�I(�\�����Rqw^ZwC�?����"Qh��
;\tJ��X��ėr � 9���82|��tH�` l|�G�@5�ӛм>�~��M�ư�Ȝ�1�|R�m�<r W�h��@gv��_&��D��<�T珲&6C��4�<�����$,REP9[�ǩ�pU)�����qir�1�R'ϖ�B6X�33-�W�����	X� ���cŞ�jjpŀ��P�;�&���Am[�xU��0SֹhƳa��e��f��oC:�t� 3��	�6��pY�7.���f'YV']5c%K�1���L5���р�D�Ɏ�p���L�ŗf����~8�[�h86��"d�-<��TJu��]ӈ���(��� eS`�6�TJog��Ue�:�p��kd̰�V��6Q���������0��ք��U��V��Ӭ��&M���g��~�OT����\y�g�S���6}U2���Y T5���:��m�|���ynp��}�l��������&��o���KQ�K|��Ͼ�D��I�#>a;z�~0,:��N���g)�u�)uq��N�o��ύK�)pP,��2qK˓[�)2P����̬i��أS���   �������C��j��*��92l�O�
���47 ���O��'�	�+Rʷ,Ъ���*.�i�=��%��H��<9sk�?5��������@�m�����t9Sj��ѻy��(���E���)�}<W�8If�#.��������uD�,�8���1'����29��B����3 f�J�e�o�e��0H�3��d��
�#��o���B�����'gJ�n"�#�@�Q��C,i䲮QȒ��D��?5�חXѓ���soy�-B�](6>!�G�^Y��-�rb]�t��NF��Rs㴆��#C?�G0�L$s6�Y���*�(��T�́�d�n�u���̮=���g�8�����}�Z�����[���<�T����sZ���a��|�"F{��)����Ѻ4a�op�݇~o[T9PwlF<wIa�]?Ԛ�XM��p��]%����kP�%��^�Sm=���5�g҄�I*S�AHώ#I9��Y9��||�W�@*�3o�s�u�J���J:�*QV�FMy+���L�@,K}�66�G��#����	�2.d��@W㠨!G��hNks}O����("cbZ^�&�k�q��W�=Jz�2�[�:@���͏i��v~{Y[s���3A[WŊZ�ACɼ�?q@�ŀ�;Q����� g�X��5���v&GUw��"��w�ӛ$�q��b�Tz�-Ջ��=\���=փ�<"�����9�����j�G���}��.�͒;�x��e�p|��f�_Ø�s�:d�|�i�˽e}4��;�64A��D#�1Q�P#��h���'��H��|N�o���Li�E��-�����$E��=��]@�����[�S�B�E���3��ݫHڳ{�d�6a�$��v�Ԛ��c��̻�,19$ @X2��Ur���]Ǹ����Y�\e��?x�u�I
}����2\��o��f�Ѭ�[sFI��\�uZ��7����{���UT�;��R���r�9�*��	 v��~�T����#c`{-��F��~V��Є�@/!ՅRh^��:
�F��4j�%���Pds��WU�`[`{���4#�g�>?N������{��vZ|��ɧC�R�g.Y�v�x�
�=y4�s�m*�6�zh^A7���a�A�Y{7��q3�$��>��u;c#���d� Oen���ϴ�/�`��^~����(*�����C�6ŀ��7vz9�i:�)*�B�c����ZbǆDӬȃ�-Ӧ ��K��![��sA�fxkOt�����#��c▃�&CJ���^��,'au��.&�'8����B�
v��c�X̉�v6��i�]Nvv�݂��V��Vf�JH�B��)dB3m�d�h��YBM�DfC�-5��O+��M�Evp\��0qh��QK�K���./��軳*a L>0mg�z
+?����g�o`CN*b$-o<��z2�
�S�$��7�A�"���hfbOo�a�������o<��Я!C�$~sa�k��GJb�+7(n�j++Z�_�D�t�%�J�{��&LZK�*�!ss�:]��Z_4�*6<�/M����@6�1�o�V���d�v��2"�<��nd=!*��V�����kt��ZD�0��gto!� Y����yK�00.��ouo[�-�擸Щ0H��;"rO�M���.���$���4e����V��a!���򽣏Z<7PY���N)\�(��?*z�����$��9�1����<�C�����U��`�y���$/�^*��A�h�[��}����H�-h�$H�t`�H}c�Ϲj�^6�7$t���G�ڰ�J.�U)��B���'�& ��'�?���r=@Ӯ�5�m��z$��Q/j���>�n��+0�%N	���Г��0�o���^��A�}j}�s^6� 倔7���܉K�:2�o;JP�'�� �r��A���їF��
�o����C��i�3EǍ�/�������9�&z��]�gG*y��c������k�µ�>E�\)��um�e�XS�be~h�i.6��W�>g�9AN�f�ܘ�!^t+��B��a��$�?�oF=�O�p���*�mh��F��N�@:�= �K#}3�z����oH.�/�FE���q��Yh�g����Wz�<s;m��vK���ʡ�UPG���8�,�����1V��鐈w���PI��~�R��}�3c���l�(��7�@γ�I�l4���"���_T}7�YJ{h��C���K�K���x9��5�z�w����eH����%��T��L%�d��Z����P��M�z�H��?��2��$� �H����a�0F�����S�Ί�'N�܍%ɍ�@*�c�G��z���k�,\�����k�=�<M�^.�|s)��K]X/E�:}�=�rrBW��ڶ`5���_1H$����5�޲��aJL#C�a�x�S�v%����/�����N� �]����L�p�N�o��JNߌf�õu%8�}�U�� NnY����f�Y	9���Th�8�s��3ñ*��'�<�����4<���yb%��&�a�p�ߓmc?�X�VI�"��~@C"}{.%��̒�a�N ����a��Q%xtI���� �������+�I��du&���B<� 
�����X��:N��4c�vkW��8�>��l�x�+�?]yb����X�H�S�ݟ8����{�fպJ��)'_U~iS����:��z(�P��|�Dڡ����a����{�F�KN
a��Suu��z�=  �y�忖�`^�!���,�Bl6&g�-�V�E���5'��� �������е��sH"#�*��J��ͭ��x�j&����I�8�D�^���J�8V�!k���: [Gp�r�A�'h�0΁rJ4?.'a��:��c��"�CShu��+.E��kjs^�����3Re�Q-�4-7�C�f���iʠ�a`�X8A;MY|�'}�0��u�_�S05�>~��,��)3/Ho#���V�Hǘn���3i��Xai=�/0(�W��>qSFFūAM}4d�L;�0Gs�V��I��3���u��T� ܖ`�Ɣ�+��L��
��m�U�!��ޝq�()��ߑ��O�O��iliV�����elV؇�7�K��t�zO�*^�)����hB���e�D���c�9]���<]�N���R�Aꬢn3��[��1�en(>���M��J�����~S�:EF;���b�L��It
�1�]9�[���Ֆ�QlV�����P�����d1נє�Z)V��N��Y=�"����pR%��I�2}v��\�*����]���j<�D.��/$w[�O/ê�r�mR�2�xb�9�D�liQ@�/�1���D�[�o�'R^��j���5ݷ���u��6��<�����*w�F.6�@��!��F��aWXq%��gP��%�ʘ��o(��e�hj֫��@;/�h�T��q���D*�M���� ��m�v�c,��y84��V���@X�4._^���U��yo[��ۑ#�[�����??�ڠ�(t�D��c�i���=����D�PC{��x\g���(?���*�7��)Ӌ}���S�6��ֳl��/j%nS��u��w�M�(�{���'}N���M���3��$6�5�{!94/dݑM��\��A�t�c�l���t4��hŻ *T3��c��h�ėd���9CG��z&V��k=�.~M�_�J!�6��:�.��l]d�P���j������C+:� vS�R<u
n�5��QNK{F�K?��J�r~��Ť�����~~�+��e�p�Ő���R��s~�?*o���L�߉/JP7��K��G�}�b�l2��2�E8\%����ad���rff�ΜQ6�cL�|h�L=Q��:��	��C4��ԴB��:�� V~0�L����}������Ʋ0���X<TM�P>%������	$΍]c��c�2�!_�tUt�☃>o�Y�i�U$�ԗ(?ɂ�@(���9�H'���'��r��<�!�<;�����0[D_f���`�g5wK�=�
�{1�B�'�]�-gu�9�X���s8�f��ʅLO�ä��C}p&���]�gf`_N}�(�0���&�f�U��7�
�uŀ�CS�v�P���h~r�P�����G�'C�Mc%L��P�p�)�+�i���L�)�{�!+�c�c���\��n�Γ%3� ֡��v� U�r��AhF��3ڟc3�c�J���a,� 1&SN��Vf��ٗ��R��6��a&j��4���A�[.�[J���f�>]��1��v#�>���/���D\���Ŕ�5 zp�(��EQ_0r�"�7)gk�\Q�`�yc	RU`%�CD�'el�M��̏�W6���m4�W�6茕���E��it��t�ՙ6Ӊ��u+�ع`�Z92�N.�������� !�k᎐���)�t�hEB�z�)$���]��R�Xf�4A�1�r�Jw��T���o/ͅ�-�X��7@��A�3���8��:B��G:�Z�(���]��%����f�h�*mBQ���X�W����l�{O�~�d�L����j��1�<Z�~���k"���v6	3�����CGr#��i&�}BE�aZϡE?��w����ٚYȜ%D�ۯN��+
N�]'�2�V!�~|+�c!hg
J��&p�,�ڽ�L'�)�n��-����I�~ii�ty��^�0��|�-�hDK��0+ǰM�VU�,�Y�PP2�J��z �96C���9�|�|q]l����*��S��E}�i���O��+�!��ލHx��=Tm^}ފw�x��/�24�f��P���6�Kf��(�,Vz��r�A k٪�%۝po��rug*��+k��c�V�8�A!�f�j�%�t[4�����EƁ1  ���'R��c�&�&(�SCŰs@۸�!Mh3r�/�-
�6���W�|T�|k��>��_�J�>E˃�1E�$e��N��pB$�͓���"��_�L@���� -k�=U�����ϯ�ϸ�d,+�n�S`����ݕY-/�f���W�܍;LV0!#���>#3L�����6��H�L�\B��M?Ω?�Y�%��ҚФJ��ۏ��_��.���%?�TP��p::�b�c� �H��_9�����(�½�'FKL�  v�2�,��H�vđ�0�Yb@ p�.��#m�q����V�� �\V���U_�}�?�=E������{�i��Hl����X!N%���F|@7�7�ࡤ�C3��?��鿠�v_�XTbz�]��y���_��|a3�h�g�Q:�!�S�x,��j��;ٷ$C���M�?��<
'*�.�p&��aȦ|��~ҥd���pO�� �e��[�2׈��L�*l~%zR<�9zJ����7��Q��eb�y_����%&`��D6�%��y�w�C�s͊83T�(Ҁ����!�X�N��՞���,� �T��ʌ;�z�L��n�gD��t��t~|ɚ�y>���j��2B�DN��۝_Q�� S��,�Nu�� ���{���i�R��	�Eak)Qq��H��7S�3���g.��8Uj�s_-��c��L!ʦl�6$�l�hౢ�k�ߜdw�36�[�
`��c�'Wed2��r���s����-W����{�b̟�U��B7��i�����ڰ���n��Wxp(o&�O}h]z�.G� �	���%�����P��%�1�v�d�o&>���I�5f��=s�q�>�(�aOXb���B�5��z��Ү
��w3�<e����$���k�}�$��!�E���2���&}��) ek�E?�9�Z���8��{��'����]����$+	}�����'�Ivf�B���tWhHef�ې�O`bmFx Gn����H5&�pMz	���(2ayy����_8�T�r�8�A��;��_9�����|������pG"�x۔O�d��Wfͦ��|#m�o�Q>;)�j��O��=�8���7�Ӑp0r����n;�J���yYH
-j��<�>��S_�Q�/�]�h޶�BVF27��>��G���*�n�Wa0�Q6�-�Eo�D�-��}!L|x���elL���.�Fݳ��TQY;E� �+S�`��@�ZR))��U���̪}�mT����/��Bs6��#uZw���؋&��u��i�w����c�������t�BRD'�}=�����}�i��tN��?t`���鄔}�x�ߟ�ǈ84�=�!K��\岩���U>F��2?V�Q�<�E���֊�S=�e��ѳ�Ԗ���Ao�gr���)p�#OD�GY6M� �J�k����9*-)B���"`�5�
ݤ��kt�D���  � ��U� t���ݱ�_�i��cjݥ&X�����;��P 5O��Cx����!�3�%=c��P*AE]~K p־�׵�%q���6�������[�x�rQ7o�� ���O���Ӧ�-䶔w��buU_p�1m*���&r��x\�v�;��� /�uW�|N|'	�kDm/��&c�$β[��f����4����w�%��,�=E,	�"�}΅��uC��*�
���]|C�w��_M�'s]v��`_�e?����3���?eb7a�17aE�x�V\�$�A��ս���+����xR���EZ6@S�e����S2��V�b�2�35�&|�i�#�����d`,q��Q18L�MrC^=c>�[H@�Z@?f��݆���fah��ڤȷ��^�y~��)&�DQv[Q�ܑr'��q�-��Cj�D"��e3�}���7���:[�M9�6#}�jߚ���|Ӧ�9D�F�g	��%����#������F��0���ə|nPMNQS}�׍2ۉ�(�����o��4mz�Y�K���0�:�y��ï���^�H�; ~�g�/*νz_��
��p� �ۈ��u�E���Q�ma���/�թ��x@�b
>ꐃzp07R*3(�ٔba��^��U7Wb/�F�?W���"[�������7_-�o,�@L�J�#rV��������S.�NRO樓�t-�L|;~-,�\��u�V^^���6�7�0�[�al#���1qKHn״�9<^����52X�!ԭ[� ���T��l�����O�e:A�ޡ"n��o0���
�k�'c�DJ�F�yM����0��$*1$�°���o��n�|�jJ��i��3;6y�Ӄ�]��X����_#�|slN�2tޏg����7�;���<C�����W�	%@��]���ND
��ԃ`���OQ�p��6"�7Q��B��.��߂a�	���ߖ, ��8������0e���D��y�Y����kI.���۾� ��f�>�������āeJ|��.}u�l��b�sy�K���³�-j����#�|����� *�%ܼ��q�V��V>�fin����}$o�_���;��WP�P4�b�䰚�I��֝���z,-�(����
��;�i�3s��3M]��]����̳�h]Xt91�@�еvaL�D��   � ��u� t����q��_������W�]X�v��H�x8�<�ꕀU��$�/ 0��B�]�B�lR�$܁��Y*�J)j^��n@|Є��F�v?���Y�e�iL���)�s���|���R�O�se�>9Ȝ���^a`��j��0@��1$tʏ��;�)�L���<�����i2P�:Bܯ�ip�ECt�&.���S`��E�ذ�kyI��/O���v�y��Ib,�^���Nʆ�㒯Y�y��P�!�.����>�o~�/�l����Aj���2��J]����N�mgpZ��~[�M���3~��lM�݇?k�y���a�G@�9��,
σ�^`��7ٻI�J�}�h���`�I.����}U^ʀ5�%��I'>�|��%{�2C�ț�d9��ө�s�z�qн����η���ߚ�YU�}I��q%�Fg��#0�?�)Df�5e�*$�N�a߼����������/������9��b�;�P8@��w:<X�u82u�b�F�5�]��&j,�>�D��������Ag�^ Ŧ$Q��x0�O��/�:���>��"�/����A�eT<9Ҡ��H�<�P�dζ��|m��+�_�M櫖T$,���8�̀OFc������!���|Ѽ0}2��,*��Ð3-q,�A���8�l��W����pTV�($��W��Grd��y��j�j� ���=��D�Y��|6#��<�R}	7��Z�o?� �����ˊ�t�s˒������a��L���L����#䓻�u��q���*�F���x� ��|�Sr4<�~�o��{�?��&�κX��Bs���.�py�}t���,��=	.�@_T'�L2��1OFn5�@�UU��O-�Z�����:���pW�|�a�B��f�l6Rd�~�j�)L�,x�:4nK�T����:��� xL,�Ό�D��Q:MD��A����ĞvZ�!�2�a.ޞhͮ�Q�OTuˉ��=�������F������	��T!�Nb�*A��i'�_)ȱ��ā���.���"��@�7aĦ��rYܟ�c�ݯ��[�9Rn���y��~�	�"�&��#�mT��;$GM������Ƙj;��uY%|%�Aā[   � ��-����4�n%�:ð�����R�J���)}V��0jR1PjA#��Fg3��2Nį�����q��"���L`��/�E�O����$+��nCh�ꠏ�[!:9���p�+T�^d�g���fe������<�@yg�*Xn����1������П'ے��$�C�ґ�0��4y��;D��A�{#�	�< ����҃����s�<��Z��� 4��{y�0R�/���8���C©��[�Hd�[䄽�ҤD�*���H
�r�`bZ��xRMT2.*uUc8��&�O/�7�&/AsΧ![xΊ�њ$X�}t��dM���}�Z��W��k]�?94'��M2]@b���Ϭf�FWƅ��%v�r�O� ���F�d{��aJ�_(\�V}�H�.:�d;~�<pF�W�/��nѿ׋�!�ː��K�� �s���N��lR�E����џ�����!������1f�SOm�"���<�u�a�g��lǸ{9��]#�J���pUA���['+��d(��dx����OI��h�N��*��w���A��r�B���0ڣ@�3��Q(гqҠ�����x�m-��kl) PSN��=+��� �l��@Ǧ���`a��9KXJy��5�袿%{�Ғd�T�,*�����& �    �!���!Ĉ"0�+*�SLp@
L�7�<��\Ug���Ǜ��|�A��)�˘�%���km{�]*���h*�w������bY�!�T��|wv��2�)x��^~.��ҙ Q��n VÑk�[��Ù��̩JK�f�;�     8!��� �̬!)B
Q(&0,�IT��V�@$E ���jb���y=���U��r��TJ��r�,�Y����M��a��,�`�m�]��cUU�FP@�i~qͺV(�<3묤g��Ut!�ĵioOK �E�!e@`��A`�-V�,�x���3��[���`!���d�bb��   B�`�8��@�Ƃ��uE"�Mw�rx����L�66�] �L<���FF��&=�c�H�&J�%Ԕ���LiB�:��d)����$����	/ ��2y	\�_�"�	��T�@o��P��?��U�<��!UQyBʇ�4  !���
e�`���j,#�f��z�O�l8#k�;��sk�|�M�*P���;��䀘a���=З;�~��`��d�m��y��hXB�.Vq�KLn M�DLa�B�� ��\u[�n	�L�*�!Ɩ2W����5���r� ��O�+�^nѱ����� �&D���0 �!)����0�aD@h4, �T��5s��Y�"њԌ���gm�}� ������曂u�<�?1R���G ��5�`�§�R1������P��KN}@K�̣  �aX h9�TM�`�}_|h�Y����Il��:�~u���9ֺ�b���)<�cI$�� o�0���։*�*��ԣ--q @ �!K�L��j!)�De%�-�{�+�[����g`��#���S�������M�VF8��"պ�kESo���r��B�Qd�_��VB��	݉�e(�2�w�!�B��U����V�vR���QH K>��@}wh4	Ţ;�O�!y�����t�9TKe�@`��8!y���1a!�%0 a��r��(�?�����N��=�2?|��Q����̴�.rK�6�H	h��H#	t�T `�DI*;�Z��������;��4�-m�8�@T�KCEkd�ǃ{����r j��`�[�3��M�R)����Nk�/7Wr�|�~�� �   ��U�U   �����C��̻Q#���QT�.����0�ӥ0�X����9�^p��Jj^KH�-g\��ZǨ���x���
�zr�(���Ȁ&�Ks�K.��p�����KZ�s|Îp��I�������gG�M���K��Uʤ�ܟך��^�ST����^�L�U�ms��v�؇��/��ހ���:^]�h�Օ	Ԡ��E�b+�9�X�kx���y�������߰d
����h6�oUW��f���,�,!)�3���Cd�U�=:]���@��س%d_����#��i����$��T]k��2^���-�a�G�̩ � �⺄x�)%�{ FA�E©E�Lt ��GP����O�KT-�%�ϳ�!A���v�z&�M�Fjk{q�J��vݱ�:��z���<��J_�sZ�=���׌L8CQ��_�+{�\�h-�8��j��z�j�t��S�!��΂�O�t4�}"s��|�*6�bU�ަe�.M����]�S�h���&�c.z�,��ũ�
QvKOd=q�'��AԄ�Xa��N����`��v��p����/�
��X��7ZL у쮝�r�L�V�ܢtG����j�5~r� *��ql�5�K�����צ��Ԕhv�AZ_0\ ����7��)@��j����=	�RjU;�_����tX��/�������r�!	2��JTyl�>9� �J��h��E�|6Q��U� �,~�2�]zR�ZZk��~`,Z�j�ڟ������q�lT���%���B4ڻ8Dl��`k��$�&4�G�p��Yc&�@D�5�{�8�����/&xn�1rX���V2�y(�-���,�$��_jր^�>E��X��l*�% �ew���Ba�Rp�O�����64�ʉ�A�'�w��Th�:���]��"��M��2R�#��h
8����jKǳ���TG��E*��|ԡ��'�;���
{��2"�JlE��$I���?������7�E��������F����h�sW�+@hf��q.L��0U� �v����������z���K�0�x�L6��Ea�YTݞN&�{���v���|�"F��(���Yz04R/U������U[Ӆ+f��P#����z��}���u#?�S찑��bN9o81z\ꈾե7ĩ�F��pt�QX�6�U�؍8)�<빱�'y���u��̿��m��s+��K6Z��%୰m���|��{h;��0	ګja�M���Q�	���7��BX�oͧ��wB�>��d�t,��-�M󙧸<�F�����J�KE�^Ϥ��"Ұ���smI�ʡ��D�4�gx��4b%&tFy�����2�~/�X��\8�5Ol4�>����}��N�!�t�B�A���@��F��C�Ww&ɳ͛u�
Eg��mrϒ\��������dO�e�+ba�o���6<t�$��~�������p/���{��,Bp����}`D]��ky�2������ʳ|y��D6N�󂀗Ԏ��w��=�1=W�^'s��=4�S%��Κi�~���C�2����7S�&���x�p���j��o*d�a�{��;��(ʖ�q�������BJ�A%���9���������&2���ڊ�ܹk�7)��k k�ɪ�L��(>�<.y��	ui.��teUrmȯ�@���pc�Pkh�hQh	�L�3�`"�9W]��y��V�a�O����\����-��A*:"������H�K��WL MKEc1gK/�����6�s}^8H�ȕ��f��z���
=���[����f�m��l,�T�G�}����?���JS�vS1�i��i�[��Y��X�!6/=��w�RmM� ���?�Ү1Y�El��Z�.��<��N4��L������hR�g(x����z��!G�g�z�v4��ױ�:�{�S�U���S�o�F/���$S�p���v�