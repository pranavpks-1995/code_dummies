�wf�w��@'@�S�&�/�i����ϩ�Y�h⾧�K�LJ�Y3[=A������-��BC(�I���;~~H��b����4�0��%Ԃv~h �&��`{�>�pH�Z)��,P��m�(�m0p؆SVX�g��P{O^�Z�{�Ū�z��E��;|R(|_��70���d������G_��-s�c����6i�z�*Js-y�����޺
Y� ����������d6�(���A,j�������P*�T!���^� ����J����\K�oKs�6��l���ߵη����Q�*�v1�c-�. YX=�v�/LBaf-|5�-���1�2��!�s��ٖE���5����x燅���z�ud�2�� �iV&Gz�^���0V=�0X�6$;<�&R�a�p��唣�H��e�L�w�ǲ�g�U �*;fQAӅ쿗��g&��S�!F���QvTO��:;Q}�x��*Lc�j14Gg$�3�MPͯ�>����q����u��%&�ƫ(f�z��ΐW/ ����lV����L�<n�i)�����S\ ���x�6	՘�p�6-� T;+~f�NZI����{�R�7X ����o�a���:(E��nG�\�p�a����mݞ
ê����I���
���ӪU� ��/c��de�{��M^�'�Y"�6�T�Y��뻼(�$ZR�=%4��-mg���8�yk�L�g7���bX]��k�Zk��m3+���Qa��4Dd/�����#��`�)�f��&1Gv%�b$i|���> ��8�s���1-�/t��}�w�Q����up��Å��x:���agK.�^�w
K(������3f"@��Z��q(�ݎ�x��$�y��O K�^��O�qρ&:�^����^�/�>�ytqc���P�����s�7(w��>9ބ�XM��I;-+I� ��x4m_Su]��9?u����/��
&뭠ű�Ko���F�^��#0�W���\�hjV93�a��N�Q��y��V2R͈�l�2`�����q�j{*�Yįm��:�'6������Y�z 6�:leh<�ozz��>�R7h�����)$1A��9N�'�U�a]�t9�������6}ENV ��RqC�'�S��TdJ�:�51��Tp
�n)�?SJ�������y����	�LT����r�Q����zm�xG��w�����Eͯ�����$�������pM���<������{��X��'ǘ��*�R���;���I�|�K�&�sQ�sKy�m��~��(���	��%�2��I�g���v_�H2��sT�
 ���� `�]�h���H� �j�-��~�Tק���t�<�ܯx��A��D��>�qٲ�b7��=ɳxAO�9#��D�+ h�(2a
����H�̞�`%s��,�����-������5�Fg92��r�|.x~�%D[Q	4_�X�WQ�i�Em{7|EN!t�O���Z �^ahXPL�i^�P��2�Y(�2êͦ�Q4N������pl�2�TRkG�a/��ȟt�����ג�����}��<x����� :7���8�q����BNW��&n3I�v؃���*���������!Zyk�.m�	ҩ�e����Ɗ�Vb8���x8 }�3c�,)�9����5֞���j�N�9��\��u�Yf���r��9�i���T�N�
��3���������:��Ӟ�'���K(k�m��A.��Sb�+��S�䩢9���&�YW���	�/Lp/\K�kzg<+��
 �Q�FX���}Jٯ�:��������M9�V����f�^�fe�˴�ܒ�[�Ydk�K�W����9v��P�ɫ4��&Њ��kB7��@�2)�%�,��H}ߡI60{^�^��@_�Ҿ����B�ᏹJX�Φ�va1re��¼�/�����Bv�[���4Sl#׎�b�;0��v�^�������56PC�ă�Ĥ����2�nt���]��$���iV���^�>f�������Q����w��f�U��|�������?�1�W��2�+t��N�	2S@��ҿJ���2OP�wo}t�¿.�(�;A!��삿��r���0��W��}+f��M=uSS�$^��H�yaz�0&�¨ų�w_��9s[`)�ܯ�i���Ę>K&���C������5h�w:�_C��"�9��> E�S�Y
����k�:��A9���ϨrM3� ���xYZ�ͮ��F�{����͠Y���������)X���k��L)�0%��珥X	k4�I�8[�8Q�t��W��␽�ף�����?�g<��es����(��X��yH��G�T3%J�� ���~���M�E�w�������V����Z�_���m���&i�94�5��9h��d������OheB׏��b���Q�5�Bix#5͝~�E��� 	r���vy'"�Rr����ff��X���P0l�T]��6�7���[����Og���em�[�~7C<���*�J?���
)��5��� w�T�yE>��a�ZN<����#�O�����LU�FF��c�8��KX�Vf���]&���ĩ�\�Y��U)����T���\=��t\'i �����C��=�,�*�}�NP&���G��r.{�\��SoVI����h���e�\3�>���y��Gz��T�"�H���+b��Q&is0(�,㐮L�nۉ��_H`r���,�wS]�\�qYT�lN����6bR��΢!���f�Zň"���{�U�N��@�)%��7)�d���:Ei�+<����ʘ����Q6����upn?!&��uU���ߙ2�wq)����c�ML��w>]���g�[�[y�����r���/�����X�Q����Uy_萛_8�xA*nX���{vΗ�u7����VV���ʑ�!c*y��RZ?kZ��כ�(}ŉ�M�(>�F�7lJN
dT�ϧ�Q���祿ȗ�*�g�Ls־�O���ŜKl����(	������V�W2�[�`��Է�ہڑ�8~T��2c��L�A�|l�Fs��l�#%<�R�7j�n��P��P�y��$)�;�3P���5��v*ra���U�@%;��Q�U
�*�Z8����2!��G^���eao������gr �E��;��P�{�?ޑ���p=�Q@ơd<��#$�̏wZ���a�`�Xp�T�{};�x�ɽ������|l��H����$��'~��MQ6/�g���b�R���c�nuN1�6E���d5}OB!È�o-�"�8�Ok|,I��)�=��u��'�j��En��<��I�����E�f$��!�.�a�|����|T���������Y	É�Y.�KI'l
�҅}⧟(�����}x"'�<����j�a8}���Ըg��c���)^�7�C��g��]L^�G���=��\ �,!�d���?<�IЬXݳ��f^)G�u	v���2���.����FV���p�;kZ�g��F��p��z�fH���4�d<�3 �-�k%q[H�uژ�����
�ib�j�6!��b��_6�So���}Fc�U�S� ��w�E�qD��l���箭���a,�2��sVk���9�<۬L�n]�����w�����7k+����)�4 ���s� 
���W��i��aK���������zP� R��:��C���w�N��{���P�u���J�x�@�-�� W\y�i�%��L��k��+�CO޼���̉/�ƽ���Bk�DDq��5g���`�̸�H�8(*2�	���s�E� ��%f���ׂ��V�,�<�}����6@�]� �*B���3ZEFs[���[O�V�Ps��7��玏�S��L��>��L�����^�=�F/͆} 0���+cNo�����6����k�dcs3v���k��\׹b���^p6�q��1�Oj�x���;#��fΉ89�[G�z�e}��gr~�~;��m������I˚���f�G���R��)�tx��CGYT�40;� �,N��u�/�2��>F���-����b'h��+t�� >�J��|���4���&M��o�Bs,H	�5��W��`r�5%`�̆8+R:��}3�z+w��;ea������x5�c �>ź#묽aH�盆�.����t��.�C�<��ex�QW�Li�$�c�Ϩo�
��}�N�h����:����-�r47��+<�2:c}'���s�y�Pn_M>zg�Ml�
X�fBKо�\9`W��0Z�{/]���sm+�R1��(�/�\}�F!�C�V7���b�Cr�]�"6�#K:�)w)��gsf�Łdt[^��?R��A�~a3������9����v���t00��=�ըk+���.i�M˄��X�+���=���&��E��y��������_%�
���|a�E��b��?@%,�es�����\�ʵ՗z`����V߄Uy��RX���[!$5jkH��H�G�ض2@Oʒ�@��pJ4�z!
��*����=ټu- �V���T����z���}���[��kk;%V�؎V���Ƕ箃m#���-��Tv囍1���E�	&j`g�g��>�r��ث��d���mw<kkݾ�1���6�B" �i���a"�T���S�eق�0�.�x�_��'Y�Mh��J��  
��B%R��c�X2[|�B��0!K��"a��1��ץ�Dr�O��9g�^�����	^��d ޫ��D��\�N�}ھ�7SY��,ܭ~���y��ݚ���C�2p�=7���Xi�^���ot�i�2�iS���&��fn��y�¶h�ύ��w���BZ��#�X�5��wL�~�mU�E��J�/�U4Ιŏ��CF@�^k���±��1e���J@�ovP���^F�G0�Ž��s��Y��=s%�	٠'�2�o�cR;�"��A��KO�|Mf�Q��LC�E\8��~��-��/��94�^L���<���t�<"��/W,���<G�:���7�4<f�Z����� m��� �c$�p*�V�f�C����A~A���I"o^�v��#dd�ڐ�h����x;@��Xu�Q�����Ajw���>���<��wW�*�U����h?Eܱ��w{7�S=�_�z���4w�j�@�/1l���s�����W�*�}!��E!N���([_o^�(m7���l"~]W�Z?�b��9Ra<;����s��9�TO���,�a#X\�m��VBm���4�v7��	�DL����E���<�kM����hu��F�.�Uu�dsQ7-d �+��X
�?p�I��0�b �#��b�#�Ҿ��Z�a�*^��C���隦$;����
d ǌR� ,����6�"]�1���� A�;�.Ո�@X��f�z�3�.�2ho.�d:�|+/fP����֖23ēcۍ�w�m��I�`���/��ƺ���@�z�	D�G6�m��z��%�}E��'3��[2��,Z�a|n��#�#-�M����:F✞k0� �6���L���RT�� ��ф.��;ͺU��<�g �S�pi���|���J�5�������c��ԍ�冀߿��6gWJo���gE'��������^,^�M��[D�i�p�`�Ri'o4�-j+#�����2�+��.��QW�
Z�4�ߡZy���g$ �E��&߹�k��A�7ӏ1-�u�H��>p�����+�tO�o��ش�3�&���	��&>�k�U��J�dTRL��۔����^b}��M�	�CX��V�cFH|W�����[��&�N=���w���"�	�ѹ6�c���r�G��+�܄F}LbM�y?�r(?����X/��l���:���o�>���v�����g=�k�22�pЋ��qUFp�/��x���	3��ь~�<�T�������ѭm�����K@b,:�baK��h�sY���|��L }�-�+��O&��7�L��J}��0��8����H�t]�������(�����U�y���ƹg�{�/���i%{�К���j,�,T+���js��KU&��\e���}�ف��p���-��.~k��s�M*��d���l���U,H�