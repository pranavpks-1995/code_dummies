?D��M�@���{��d�0�y��/�>�Z�����@�#��$ikcJd����0PIҷ���]f� NA�͖�����|�U�u6j�3���X�E.	§�c�t�Q���%3���/eq��������5%ׯ�-K�q���p"�6��9�BJ����Aذ,F��d⁣���f���'��gT[����4[r��R�q(m�t�6�+R�t3{S�%��r&��}A&E����^��þ�f�ܞd̆6`d��va�7g�帕益�umy��f:v��:���
�=���t
Ա�S��}l�ֳ;Ɯ��+���P���nW>N���U�\f�B�f6��t�5R�]~à0ܽ�^x׆B>4�;z��pkS'�&T{�:�+��Hu�mqpC$,�@�nM��Ha�.�/J(TL]KL�����V6�fȕ^>��,�{? s�q�l?�èɘ
*F�*��i�F�S�dO���mݥ���x�! �/e�E
�ii��d�T�ع��O���R	]fh�\I#�>V�ꉻM������#�3Y�LDЩ\�[��S*�`@b?f襈�z�0�i�A]Y[�̗�Vv=l�עզi兩A�M�n����)X=��}�:�q�Z߬�}��'k������.�@��$aGiTI������m��l���p��gأ3���s��,�����X��ʝ���31�|�qz�7��uE�O�
T}D��c��?��{Zck�C��A�W�h��H��c���s�ұ��\�ٹg�9��Ά5ڗ�_�6�4��d���)i�W>�����Ԇ�,�~Dw�d;���JR�����>��)+�Τ����wp��$��E�
�d'���:���K�p��3M�JUR��ܸ��<tW��|��>�{r�h�m�vA���u!g��m�7�0jgL�H��1ہ�>�_�+�����}��pD:[c���;�'�`R�̒=��r��.V��1�%;$��y=(Aa�1�ڧ�'ǏI/�ݢ������hoCZ^�2�&�s����vw ��:q��Ω9��!�i����� �m}�>tu��B��B��疬�X�h/�56��˔怙� �hc�\��X��tޟy����_ ���|г�[� ��N
\^5T�p3�n%�?Jj�ѨE��Б�-l̐�A�)�m�S����a��ka�������E�!� "�A�����UnҥA�lxt���lV����JK��=�rIq3��z+��4��,m���^�H�-�=�2'uti�0�ź��5���@鎜�QIT�� n�֛��?[��ɭk�x�D0�n�K�"j]��dZ�:�B9X)�mE�$6ګԇ$�$���}��4��ʬא)���;��#�̳d��V�].^��c���IC��W\�03���N���_��3J�������.4;.:f;�Ύ{�*:��'�$� �����R���`4��=ҩ̿�%
���G߿ 5��d��pL�n\c51[�h	qXؠ���"n,�V�@՗���0�8T�E:b���^������e�YhnX���m��W5GI��ʆ�)aė!�`bI�d0���#�;`��;,@�F%�Bۧi6,�c�zBQє[�/���~h�"5�<�p�{f�q�q�}��ƺl�	t8�����>�ϭ��M��;ŻU�άŖGG�|t5����,��f��u�ꩣ���vJ˶���9D.��N��T�E�3�8K��G��e}��n(J�K��C*/0bk"@�`�]�~ޭ�s�؅��;j�6W@¨$ُ�C���]�T��? ;!�>��&�]:13ޣ�Ȭz��?8�����f�3Ń,2��8LD�k��	&�ØDCE�Zi�UuE|&����M<@宔H�8;��I�o�|j6/�x�Q�ᒁ��n&�8�1�
h�����X���i��\״:Ώ�kȜ�e�>�)��7Al���;�h�ŉd]�,х�D�İ�F�E�y�����t��������E�ĕ�JV_E��i��D^��B�dK���GK�;��sK�J2�$�|z>�y���0L{����*�zB�m�v2��rx'��_U�=��f��pGV�ЊN㞘+�0]q�6�M}��H�4��+��C���=�yYh�1�S�09�V;����'Ǫsź�n�4���H����/�����%��o`�r���`��k	��������\�~x�a��A�j*Yk���J��������0=F�<��La�W���\�)�W�Lk�\  c��%RW�c���R��6�]�П�X��2>3���B,a����SLd��#XBF�O��@�RK��_ղ,��eO�u6D�qU�D\IJ�V5@�r���MV%�Pև��.4KS��>�aK��h2���Y��p�<�ܹc,��g~��!#&���v�x��Lz��b�@�y���ZcX�Ê��53��� ��,(�X�q��^x�؏���q�����e	�1�n��O����e�����
��\ÑU@���fJ�)�-rD����L����8�Ə�%�ެߵ�s�x?����-�Qϯqg_]��a���j-bqƩ9I9�AmP�Z��Ea��_kf6�f�R�5����'�y(�Ae̙�L���ٿArb$"�L\�P�{*� �
�
,���c�D6�2f��H%3��� k��ǎk�b��T{���P�UC���[�y_��z8@z�p�p[��Sx��4��'R��{��&��nH��萘� ƲU�W�H�a���qa`��yу[���Y����-��]�����p�p�c�xM=i�.{؎(�)���5��-�=��?,&O6�w��6�{��vz��g$��?քXA����]sAu�M�!0'����wT��9N:w�%����Qs���v&�	��W�b��p���"�8%�N�鷞{��	�=��fϞ5r�œ��\p*��D���\�Q��O���Ɨݥ�,6�	8u�U����e�oS��E����]�Z5׶-3Mw�_����hZ��C��:���o\kaf+z8��Y�%ڳ	񶜩�!5� �ը��v���b@� �]��Y�|F��+ت�nX&� 6ճ�fHB]n��X5�A�L�uuGŀ�+�;z�0��-_;d�4|��I��˪l���֯!�{�Q]qxB�=�9w�jp���o��U�����6jpm<yt�Y�js�K%�s��� `3�
�K���C�)�1s3��<�4�oQ�  %I���{x+P��c:x��GI�\g7�n!`K^7���D1Ћ�M�
v��c�c�Q��y'b)9����I�m&��{��'�jr�V�F���I�V��P��LhL�U�8W�x#=~�Yݸ�^�ԇ1���4�ijMh&�%��%2��vD�?ȊW��N��������Y	�Pa���
;��,-|O�
��/6�w^�{�C�UvM��{����� �R~CS.�������=6_G�}9ʚ.0L�{?9[�R�hzR��0iSS���/lN�NE<�W,yt��N�;0/�3idS�T��W�:�T��zP����2A�����4�r"}���� �}��X_�?���0�8�9v9_D�[��w���Q���9�����'v�͵z��̻����Em>�6�����2���8�2M�߼�l�b^ �+�#�z�|Zbؑj�"��D�IZ��xl���R�ۅXm�.!��U�W�u���X�5��&�<�&s���2D��I]-���)U[��ȓ��!h��_�d�|;W2��G尮Fc�}���&��
��4t�V�k��uy��`E���޿��R��A���}�-���.{���nS����V�Ɔ/�"��h���š�A��o���[Yf�|��f�;� ��x��T�`��Bi�_~�0z�!J����M�?^+6�m2�7'��E¾�H���� ��i�C��9�rr��v�~��ll�H�t1䐡��*�Hp�/�(������q�:���;�s�3f�]P� ^���a���"3
�i�]���5KA�}Z��~�D�v�Vp����S硈��~:�C�<{��{r��Ya�>���Z���q(S�|i���'������KV��:��)���@L���d�OP���m��o��r軁n?� ��� ��=�g1��ܟ�T�R�(�,�Rl�6�f`�t�|�*��C��7��%k�v���M�.��Cp�C�9�R�n���o��{Js��T��3��˳�e~ز:�j� ��bdNj%�q9��2���Cm]�<�{�]WP�����fdC���g�]�I
�����2y�V��:����2��j��</+{\��j�ܞ/�� l\!��*0p�g�����J��F���������*���6'�A1;�
u��Il�j��w�1��8���DA@,cr1>���Sy{�F�A�Z:�Va�X���W�a��wc�Tm|���\��mS�0�^�r��R�h�|�%¾�^��=+�Vh]���]ve��cÂ�T��U^���y���J����L ��������)
�֨X��P8�N�y��n*L4V$GW�0R*5����cD�ᨶ�?���J�8g*>�-Z���,�(����b�$@�S�J��rB�ƚF�GP�ё!��+\h&���U�6R�wΨ����+���FPp������q3��"˨�-�ӊWhi��EOH5p�٫�����s��7v�drޡ`�Կ�P��z�-q���#��E�F���t�|Jzti��6H��o��G;xZ�)�-Ar��ҕ��`�����Q�;�(�8,���W���q@)Daɏx�yt����Ls�(�}I������T�j"H��{��Yy�o���|>�Mq�T�kx.җO�`7c��pL��6��W��Xӓ�m�{�t(T`�������i<���`���NM���Izs�߮�/�wW���	����A ��&����ٵ	��5�8�w�W�L�M�6�E sM��9���}DZN)��F�����*~d�ϡg=�f��!l�]~�����m G���ӂr!YXKvJ~om��롟m;�+��7w˽���u��W��j5�v�`R��JLBR�F���~����'���=��9�b�2FI�|Yk&WV��_�O��BG����1&d7wZn����=2�6Թr����N�I�"@��7܄����*����ib���
�g�|jiꚮ~.�.CFOy��c�������Y|��>f��X������~Dl��ǝ�T�輵��F����t�z�uR��9�Β;�*�	\K�#�I�U��Z�9? Fhz�����њÞ����h��W�|?�%�)��v��~���㠣�)�}��h�