M��2uڼ���Jw��tr��5�Lՙ�5dO��٠aAM�z�M#�U]�^u:�K�@�}29�9����ucXN�і��*Z>9���]�8��4<��N�|̍�.@�7��3=��,�����fߡ��,�1�O�7P�^@��*8�j*�A�NCVϤ�6X�U��nUvH�.Cu�|Բ��ӂl��������!ǂ?��Ȯ6\�kA�l�UC�!W!��xo��QIS7ɒ�| s}�F B�zݫ�b�"��͘4N�i`��t_�4��T�Uyo�h�	�u�y=�0tv���
���*�����O��+qq��L����s+���5_P�W���_T�c���O�Ip8�2k���?R�x�Y�ܬ���(͸��Y,��Հ��ׇ�Z�/.8���Z��p�$�v�:#o���CX	}�lt�yb�Ke$6{hϑ��[ ��o�b�{� a�׍'�5������|�ǹ��97d^T��t�.)���/-wǮ���Fq�;�X����� :4�G�G@����.���]��>wI�3M��+�����O�	�.Bq$���z~���_���TŚB����R9�~���fܪO��zҁ��f�F�W�95w��~5�<¸>9��4�B�G�������i�2��(3�6���,)�F�]���[�L=���N����揥�Nu�{7"�+����,p$���^����(�'����ߍ@�#��s>ҏ!�Vy���TMʿ񚱾����fsI_��[�V���,����5�,5����TO�;�VM�����F٢�T�]N	\hO�km�,�N��У�`j�EGzy�K�E�%��W���
�,��L�#nN�O�������(�3�?H�4�-�u<H���cz�D�9��Ġ^SAI�c��ttv����z{�2�4��~�%A2!��UR7�1�λIL��{���rtþ����<݉�*%��[��F�d7���w�2&ԅ�ǜ��>��%��(�v,��}9Y�veU�vQ���!���^��Jj�N|4&d�|�e��tЂx�t�_���;��r.$̓�8�*ӕ���O�����\��`P��{'����صx�V�s%�|���(�շ8#u�d�؆ ۹~MWg'����r�X�������£����}�BnMb����k����S7��A��a& xAW��E�ɯǠ6<#��]L�+�W7�ɹi��E�,&f��b���y�*�Љ_L#m#:C�-#��R<��:2��'�IMq;�7l<�L�7�6���r�s�'�R9����;��V7hЁ�IGG���oMhc@���=H��