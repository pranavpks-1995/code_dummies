*�����RA.j��|��i�#|y��D1Y��� ��P��Ē#S�:>�r�}�zB[uK���X��S�j�XL�J�@���    � �B-W���Ze��������õsJQ�J�Yz���.܂��ˠg�Ơ{\s�c���7�@5U�����
����y�t	e�G���W�o����	�`�����+��]h�zҴ�*��.�@U0z�M�/bK  �$[�Dc�}R�r�v�	����K�Q��w$�i"]�r_]�2�b�T|P��0�f��N��@e��2z���J�>�@z��3�p�@Ɏx�U�\]z�F���C��EH���������!�R\Z~��`� yڱn3������&�r}b��˃9aɫ�+���M��u��V̄�G��RqY;a����,k��B�c ��'RPy�Ek���U��	�ƶ59�_�����`���b�]�[u|�!B6�;
��", �L�Ad D��i�U�
�3M0� p!�Y��I ��V�#����fs������K�f1�韃�����J�?p�~єPH��[��ѷ"�&�
�x���9 5�p�+4���pĝ5����*�� 2��S2��?o�SU*�C��f,�@�1D�}&i��|�V���u!nۚ��~�����@ !�m��?�	!�	��� e0&�=�*�c(qL�Pz�k��.���	��O��wN�!1K0V���i2��p!U"��5�  Y�@��|1��J�d(�\~�����8��]|&v����d���	X@\��a ��6ƺ�� �Z��<j�\�3V` �!�H���6 �˺ٰ�F�t��=c|��q��)������|!q�bb��te&9^!Af�!�p�kK�E�D�9p�L�q�AJ����@l ��_V�>/��m�����ۙ^����넂�.�w 8NR�4Qi��Nҋ�P���[���2�T���嵨��(�\mG��s�]�*� �!�R�,��z;`:Z��{,��m��ž��(t��Ag� �c=;��n ԫME���@;P�*�$�$SMֹ$Ea��҅:@h8 �iҶ��C��;d�=��v�WZ�X�;�x���Z�y�
��U}TK�ʄf2��	�Y���)�T�+m���y���wr�I  �!��H�,
� Y�	8�$�A�b�CGL���UAQml�p���e�B�8��~����k�!L���	�P��q��~��Aj� �H	B� �
�`PEJ