~���34��+P������Ǐ*Ҵ	4���q>񅬪�������0�sl���I=�ͪ�H/�1h��[ ��X?v]�������)��=���aT���Ëzүd�n�#�*1b�����������P�L��`���������UV�Z蘏Y���֥�¨oG��l��Bj3J��гҁ��a�#�Y�̧��[sK���Q�yL� �Q� ��!�M28�p��= m�*o�-
��~2  �6������[�1b�"n-�����~�h�����C�����{!d�t�b���I�Ȏ���G��e/����� ��5{�k�#k�qǳ�������V���7_���K�}�'+�jz�<,�~����皓ׁ��1��ڞ�D�%>{c��}��:=+�T�K!���@����Va�N��eh2E�XT�&�i��x%�����W���L^Yi��۞kz[���\�HQݥ:j����m�V��\\"��R�)@�Sk��"�����d���E�s�������p�윷i�ǈ�ʊa:=a�D�4���8��vA���Ӣ4d$^�ܗA��3=u,OWh���9EI��
=e�/��u��в�pV����.�Qk��C3<p���71�j�'A�A���  ��'R��c���Y/�����o��"�3�&̃�6�>��vF���nU���9�=q'��F��ҙnH�w�p3�P]�o�L��:����%	(&�E���}�!�8w\j�w�ZeD.@�"���U֞��Z}Y��5b����2}����y]�ۂ�
�ɷO�B/��q����@��	��ֺ��Od��+����&�P$O+n���:�h@7Ou��
����V�kˊ�>7W\X�hZݎ��%�N���k��_��=礭���R�!��G"��\��p�]�ۓ��)�c/K�
NU���9�@zty#O`�y���[��͇n�G�dy�7U=���=w�^�~���gM��B��n�ְ���2ې
�N��d���ҟ�b�1<���Qs���a��A��h  } ���U�y�U+*h���@�lX(+� s"�u�.�.)Z!)�3z��i�� �q�������j)�*s.����.=Z71�Q'��y���ȏ�5���7��^���y!
��V�ciw��Y�7"�`�V� 䑣��5��>>�de݈����n��n��,9�p�602����S{>i�ߟ��|�Y��W]�ɗ�v��I��P�ܦO��F�9�qȴx��B;�Ƹ��EŸ@��Z�F��ƹ�yvX;�5D/��(I�(56V�E��t�ZZG�<ec�P��Ld5�� �쬺������p"������T�P@`>V�$�ΈjO�u��j������fX�е�?��9�ܪk(>HBq/�&̓��p�Ai��   a ���u�xk�"p��@�_A!����h��^�h��ϱQ�����T<]Yn�F�D�j��vR��	��n��$wT�W����ߔ�ns�?��,
�y���.�Vה^�S�pF��<������/�$�Ɉ�Zo���=c�$j���d�.��z�{�'\�Hc��[�}��}���˅GwN�m�Hf��2������`	\�P��B�Ml�tw5ސi�a�����p� j��NK���Tى�A�#ۉ����<���qo��i�ْ�v�ig��ٻ+�p�p�;�i��U�eR������ُ�	�x�����)r@	 ݕ��-HX2��n0�V"&���K����4��@݁�    � �"-����՝s�ԭȀs�7F��0Z�r*�-�r�:�ǧ��m�����U�*=MӒ:j�'�1��߁p��ׯɓ}��I�/F
��PA�[��>�� 4�g�b^�8��ń�!huR̗�ӊ�.��F:	�G�Y���z$�o��u0,���Bo�/�_���"�/R&)
�}�t���c�t�%C�ի 2�N��Q}4����+Gȳg��@���!���A���hV
!YYyaK���oSK`+1ʒ�+����D������t�V���y
�"�ܥ^�@û�"�n�a�ⷾ\?"���Ss7hѡvW�>���Y&�$�����Jp�[��L@�CӠ�sm���q��ݼM�� [X��Ɣ�w��C�Fu��   C�u!���T� Pg�  �  P_*�l\��D`ǘuG�r7�G�lQ�8��ˊ�$a��8�Yk����D�'�Q9�/f�?碊�Hۉ����n��*�RXw�k��k�ѹ�-�o[LC����s�N�z���i�W��o�"�iNɥ��A��&L���+5S���K��.[qz`wʜwŌ��U.sS�a�q�bs҇?������i �ט �&@%�th"��'q�/��A����z�^bi�c.��0�ί{�b{	p�E�]x�~�ߝ)&�4O��M����o���3���5��3�����_bD��ݑc����uvщ�j^Z���{��Y��x��c[Q��������*C��+�/�P�j5;���_�2`.��ßt8�*�Ki}n�	iR���Bx��'ءp[k���bp�I�;�?L� o h ��uM��26�����ݬY�Q\�aޛ��t�*�0��W�i�߸���a
}&��ͅ_��ʹ��3��5����	���u��
���Bj��pȵH6���`��"���)e{b�����T6A�a�(
�O��b�6g��NB/�F�ٚ0���3����Z��b���N���B�8���͕FMȀ�m���\k5;�X��ιO�R��P�k//�¡��Cc�B*3�+Rw4�"�s�:�D�s]�V��U4������3��Qc����\	�6�k�ǖ� ��ȣ����~�37�ϷǍ�E��2n��d�ư��ܜ
����E��/�_K�獱E��s�W>�I�G��N����w���F�⻢�cL��X"/iZ�bRK�΀�d�y��#V�����j�Q�@+~F[&H���B�<�\)����ǯ�LaZ���0v�E@�����V�O�eU���m4�++1P�<O�̋%%1���O�c����İ�eu��l����F��Q�P�h���I#!���h	��Ku��#�RŠ�)��"#��ެ����/�^@�{$���I��"�xwK	e~a=�DʍQ�7"��˶����t���e۴����q��PЪ׉�B��.W���E����P���<�̓ނ�Q�w	ʢ��p�Y@��I3�n��8�9�Η;�~�_�./�&�#�`a�����걺�^� �e�#C"��o�W�S�Ҏ��A����X�#��g��t�ǥ���e��SD�iٚ@e��}����X�3���n��ݞx�ȕ*VyӶ �F�u�S�c��+��
�S�n᤬�M��~��]Gj�3��t%��:�&'/ ��4K��t|<c^?2��dNZG]S���Z	�	kJ�K��"P����Wô��O0]V.,�E��{��~���I@�ϱ��꟱0&����k�m�:��/8�o=����D��@��(1��[-�i�1
Ҳ���Ы��:���1�6@�j�J����g����3��"�ׂ�����j\c?�B��e� U6�f>t�B�<��L�)^3��%�a8����E8~�!�㽻��p��Ӈ�,ʀ{�yb��	2�����3�2�N�L�L\p�7҄�)�N�W"Pd����^fgU0�F�D�^���3�7�D]�r����k�=��'�iM �>�w��� V��v.s%��"�Ϊ�5���R�1��z9�h�{i���R�u�haW�☶��Ұ���+�<X��K ��7*'�>"t�4\_;�$�&�$':4VӅN��8�U�������I������~�s5��i��xS���a�0��XFo܅�A �����8��0!S>� dKM�4�2d�	����7xX�`�C[��O7�:�Oc2�*Ӕ��:1�)`�l�%iK�a���Y~�y���/�xwɐ��8��*Z�{Ɨ��o��8s�&t�	��L��a���T�L[+�r�{g�_Ȋ�ϣ���N��),[�z�Vo�z��%oO��0���;^J�g����uF��^j�Dđ}�x(^�x��������WT)�� �������)����|�V�>]�8��U;���RL��T��Փd�A�^QxQ�e��H��
I'i.�<P<�1-�����R��)"5l��9e���	-���c���h%��(i��,��֟H�y0��T7�J�.ݚ��`O�+��/D��&y�<�	�Y�h��ZW�a��U����TX}�{p������l������������ُ�%^EM�8FI�ɫ��o|@���8�(�VqᏖj��ԊEC�N}A��k�ճ�9�\bV��`$�r��m�>m��!�EG��C�޽��tP{�L�ð>|��䑲 ��ۺ-p���P�d���~&�Myh,b�a�Y�{RצԱ���F�D�r���J�w-�Ho��B6��{�;kȥn���Ŕ�W��!���5�L�l}D��f�O��\�µ̀:ʽ=�h�I/�+v`��c�Q�g�bO�/L*��7�j��;Y���6Dj�-�2J�0'��E�ۀ��Gi+1(H�g�>��������x��A�F5tjg�ق�iL �Ӏ��F�Y������eg���Z?=�{��M<:K��
�[�{����)Lm�j� � �u�v��sj�W���Bo�ڙr�!��EQq���E>�����0����
�Shn�����)��}5@����(�?���Z�j%�$�R���L�Z/M�eip�N/���������޷V��p������R�:s,hvt�F�S�ńB��+iCc��$L%	����h�&_�ā'����l$��E���a>0fΜ���@�"�1�%`f�>��˗&	|D��$$wu��E���Q�R#�ľY�eRF}�=�@�}��1�%��M�,���Z��W*`%J�~��3�Vx@ƒƅ ����Yvfŕ̍��>�IU���h��F�w�U�8S:��)���8�Omw�@�̤��'@]����[���X\,��� g�Kk��s�T�?�i�J�#��Yתʽ��/k���`y��;ѡ�B�mPr�!l7�����#�⏽��c�>7R��d��Ԧ1�조%'��@���&���;�p¯�m�����x1E��uҏ0'j,���
�d��k���<��N}�-7-[?'�l5n&���֘^͒ ؚr��7�Y�x(MB�G�c;�R5���w衚[���ש��Dà��#�0��~�~�5��d�O���j�V40���3��j�^�+�eh�Ͱ�X�����8�o���Af���3�rnN(B/̫�.���Ad.ޫ�)Կ̿J̜��ۯ�Ĝ�����u�n�.���s�G	>�N=��!�%��2�QC��ү9��?	�ϲՀ��TSN��7�e����W�u-�w�c�KS'�g�^��~"ƭ�2����!��E����1C]�Ul[C�,J���G�¯X������v�>f+u���t�ʧ�C-�p.S<���}�?������#��	 5��_����'�J�1�S{'�>�3�6x;Z��>�x�T[��b�l� ���@����y��U�z��B(��(EE�&��������->�U"�?�?8��/{">�����yܳ�ֿ�5Uōd�O|���a���[��f���Z�1�yCK�U[$
�k���`h����t	�!�!��z[�N5�e:J*��z�)��սk8%l��UQ�'#�t�@�v�2[�sm�6gB�e�+x��S5�z��"��������gj_�4������m�-�q�<��ب�'��$��ګ9O���M0*b��
^��?���W��vΥ�+5�w�b�zŠ>nc��~��6D+�'+6Ҭ�R�Je�XK�q�=C�}��NF%�t<��/pY燞�tS�;e+�����s�K.��zE�f��2b4_�8{8���ͻr����W���=�,Us%�sm����au|�)9��s|t�U��� Tt��V'�����,B9�Tv�,���������������H3w&����G"�����[�J���W�>�8����'�!`܌o������I<hQ=eF���jߌ�t3�g��@3�[��I��:���p�/�Ǆḕi#�0��A%�<ߞ�@����|���Z$�Ѿ-`���m�c'�>�����O��o�C�'w���wb�g��K� �%����j2G��z���g'
b%< 8�T��+��Eo�ǶJ8_�R��}��T�C@��V<Qش�����]c�AO�=B�L�m��.�Rpy�&���B��f;�.#��.%����-�O�[`\�ڃ�tB�����ь�Us�<
,�
k§aJ���������O4>{�-�>�(
���I�a�c6�5ğ�$T���;H�l�Wxwh,�XK�/�#��!������%�����hNK�Z�Z�bW�iL�/C����B�f���Ѻ;s�U��Blݵ�J�/k*���S�M�H�0����]:6ʠ�`����r��|���U%q28�"D����yB�!`��H�/���C�~�� �#F�c5v��|�%�51~Q������ݾ�u<H졶mŶ��_8�h��A=�w509v�|���)����$������-3Yx`�
����2Ř5�����Mym�L����Ƶ�ٍ�T��]�y�T�d\kI���>B��;��'� 