package PlotResults;
	module program (Empty);
	endmodule
endpackage