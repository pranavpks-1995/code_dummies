n�,��xݛK#�y�|��u�N��\e�����4�!@�=W�Q���ζdZyO�G������HAT4F���і20�JՁ   
��8�U��C��5��t�e_��l���Y�٩� ��n�]��)I._�AC�V��²�p�Qz�W�|�}4/%��B�v��Д�#��\imU,����`!�r-���ن�s�x�Z6�&�:%g���֫���i�ȂKg`E���㩷�x9�K��hL��鍌�"��Ol�E���wjcv�M�p�����T�CE%_:@�h:�����X�fʶ�׮�����l��(h�B��"T*s�a���T޵
5�I�F�(�� G�AR��%�^g�,Ӫ�����&D�6:�S����E��ܟ!J%$����P��WM.�P����㠫� 6��S�w彴~�Lmc����P�tխ�9IO�^�5�.�VQ����ԟ&�j�Q�%������A&�%�!�8"�7��HI���3������-^"'�񿶿qp�r����g{˖�����>p�Y�ICL��\n��!+W�˃M��1������x����!G���e~�κ��N8n�Z̡;��?�p��<mˤ����2x�fM( }2|\n+7�mt����v:���@\������2W�H� R��-ԋ��T8�>�K�.@��2U?�3H�i
({	}Y��3�_�?��x��&X���ϋI�E�/��!��*�����d�/�������5/��@�+Sx]XS`�XBߪl������^�.,g���(�12�~�P��*Db¶G ]*Hg��ח�kҋd��-�wt�z����x��#�
�]5�K	�