��[��>Z��3�6^�/{k�|�pZr���A��̔4>��&|�}���#�� �:���4���ڿ�}�Ά��(�Z,��=�0���T�H�Lm1���-2&e�<��+�E$�Y��I�oF''��ʨ�����l��+m����GrB:�$�٬hn�����niF6]8��Y��l��%K����M���I�18��)CF)2�so�_K����Z<-��uh���6������1�1�
�o��s��۪A͙���������Uq�).�t��֨x �����֬^�}{I��i���d]i%Թ%�
(�:}���`�Tf�{�0rjOo�2�۸�H\����E�����v��=���Ae��6�ͩ�Pă�<��$"��91��A��er���8���A�zub=�S�Ȗ?�#YC�V�>w�ܻ�El=�/�v'����R[����+jѡ	b#�'O�u�b�LFV��peq��7!�A`k�h���5	��H\݀�p��4�+]M�ĳb�;���u:9~1��t��_z�o�o�e�մ�LO*0�-�o
�
5��u�bi!��q��L���~�=�PK6�������Z����i��k98m�#��ؒ��W�)�x�<�Y����Y3�v��/Q���n�D��'�,s��2��������$���P�{H�4�l#2Y�x���G�v�=�m<��M�$)h���@A8���`��-�f+���Y��t{�a�u�j�dz׊A�=�Q�Z�v֎(�����0�W#�C�7̈́����=�����^��8nQQ�I/Ea�`)g�9���!n�)����·ș�J}͙g��S!�fsQ�/*��&W�iw�ǹ��&Iy�k���l� !XlBY�;�����+��:�|T�#�*�%z�X�N�V�;��J�ǯ��zx~�#xFN!������&QekCz��X7���ҽZ[�B�T�V�|� 'aMW�̻(��3m4_����[�������Q�f=�(kݺ�5��1h��#�=�sR��x��� 8&귪�ԃ�}v��
m
�B��������W�?&��)�1^�1��M�4,���
��yH�fХ������v.��`��S��G��)d,���H���  ���%Rq�����tX	�z@� ������,05�+�N�ȹ�O�W�ǈ����/>W���L�����̔�ke<�|��s%&z����1�c��+�,I��Ä��!����m�!�ٗ�1����2�+�����b��31�XN�9񒭔�]ٖ��@�>(l4�<�iG�_;���w[���<��5N�d�;(m�������� Y���I��ݫ'�f
3ݱ2Z-�|�%�E_�ǅ{B�{4#�2�N�x,�=�~�CL�9���*�.歈Y�D�rJk�]�H�^¾�Lw@/���i�C�I����,�R##B�dX)�P���n�����}���9i���)݁�� ���Gk�q4eYל����$��#�As(��ý�Hq{�T�.�&o���g9�t��%�u���\�q�I��QB
��C��D 4����Sq+4:���p�=��Y�_���qk���G�Y3���M�QT3'��e~�T�J܀�����-�o�|��T8G��d�����~a�nG��>�D��<�$9J���SL��%c\�9C�r�-S !�kRy��
.M���W[V�eG��<ф��?;��d�O�u��&�l7k��Q����U����������|�