E��-(կ���������H���$g	;"1˾��:�$Ǣc��<�,�P�� ,�o[op\�o���x�����.������,�]����0IL��^�{��zw�d9��#�%�K>C|�r����4��U�9���z�j�3۷W)����3���kmdl���H������)�؄T�uI){	@9��釜��p���*��1�#~��|%���(��d\×���(U�:A�0q7�ՌP}E:�R��C ��������V����ۉ�*��Yax3)����S�dNZV�7�����==xQ'���;* �ő/��!bke�򦻣�D��y^���gkb�[�߭��x$oͅ�A+T^0.n����"��8����w��z���z�Sh���l���:ހ�,���7�9�ϩ����\�pr�޿Q�]���ɂ��糢���EGt �+~q#��#���s夥hW��⓿L��x^�8 ����Q�D�RM��E٣�f����'��ՄyFDDՈ�[A�}ٸp润��\|�)��f�e3�ߎ������b������j� ��Y٬{M�D�~~W����D��#�S" �o��?������I���|��k��#��@yv���*��>,B����n�d���Ƒګjt+k}_�5���[⋋ڇ�*�z��- ���I\ӿ҃ن�W���w�o�Q��Y�	(o�]�L�qr �4=	V�yx�@�/�x�������.f)���BR��/1r5񴁹>+����"†��Wu��Z�ʀ��ťJ�A���^141�k>�6/�d�%݇�Z��.u,M��S�]m�SA/}>v�ׂ�(�ڸݘ+��<�M�.��E�E��?%�A:��8K��%�����64&{5>Hd�҇���>�W<e�l[t����d�����4J�8�M������<�3��

)�tx���]�?�a9 ���2>h ���ѳ�XA�H�A"!4��	J��^Rn\��`^�o��fV��E�˔rm�m�P5-R\8AyR�q����1.A!SgY��pb&�o H�Xt�I��i��=J/!Oze�1C�o�4^ ���%�B��%���I�g�1�h�,�� -'K�\&��z� -��%Ƕz*�\��1�l�Ms�:gxD]�o�z!�=���H��N��z������%�X��"��,��� ���z~f�(��p|���w���e7_ti[o��{�>1����/m��	��q���bEp+��_�����@�Gv����c
'�C%�.�D^;E,��_8>�J�r�	Bv�Sב�K����Wcr����F��ֻQ:d��n�>m�P6��V6�K�6����v���b!&��T$�%�j��Tt:�ZY�X�0��,���
�]��g֓�<����"�2�����Q>�'I.�����5  b�η��h�f���×���r���>\�G���f{�6P @���޵|M��S��NGA�F" �)�_T�|��z�Q�Z�J8�S[4a��6wbR��aX	X"�^"���ඹ�U]q���!G2���?@�ʔ�E��)��kF�6Tnz`�)��F�C�"E�/�f�|�M�<h�[�1m��}HpU54$�T��?����P�L*u���x��_4q��
&Zh"��e<K�ف A��s�;ESe�|@��_���-�Y� ��S^�T��o_~D�/ei���.9q]b�$�I:�E�<�����z�����E���~${�{����*��_xgLI�]�%��Х�N�oK�f�j<�� �J	p�?��M��ڹ�4���}����B��f8��;�������E-p��1�|0p��	d.��7��	�DŜ	�f�v�E�^�Φ�:suն�6ܔ�*`�x�n
�=qw�%?�f�e�D��5E���Y�r�lΉ �9yRyyHy���}5��J���&�@j�F>�.%�� ���bw�(�P*��;�hU���J):�`Y�>J(`o)��W�1�����Y��c�C�4��c_4Bїa�7Y�".�O�x�c �?3�G�|B��=p�j��{wj)E�"}\ x��r���r6 ��/���ڡ6�t��_����i���T�!N�c�9��œ�=��N����l�GZ����#M��e�x�?Ǿɠ\����i&/r%Z��g��V:0��4���b߆ 
#-�n������O��6���<�Vl���EK?.�U���o��jX����aj����� 'w�=��R�t-^�oY�t��,:�I�ڴ�-FS־9�5��u�	S�Z�:�1��i��[m �f�ѥ����B��B�xq!�>Wn['y|^�jTH�q���cB����2���:������:���.����B|I��e�q�����׍!��"��W����n,���Q@ms���'Ч��S��{N�}�wZW·����"���y�Q���MXقd¥�DsUǏ�/�VFZ�a���g	V�v}�������86�,�@3}��h�:]�D81�u_b|�:Iƅ-�vLE�~�E@q���a&�e�r=VA@wnT0�����*D�u��O��m�:��D�{����nS������O+j��i�"����z�eC6��dp�x����WT>�;����[f��z�B����Ez�����'�!Gپd!��.⩒ߌg��q3�֭#�Y-���78E��SKl�OD�b��Ч�tIp��ф����6$fֺT��Ė�F��
C2!���	|���w7���yy��#�,Yl��"��a�ErX>�Ԍ���9w��R9�jI	��g�c�J��Θ\tȋ�'������ƮL�@z��=�FИ�X��@��U�&
ֆB�W����C�b����&!Ϙ������0�`T��d� ����
c~5����`)X�L��KV���]b�2J��K'~���Z�r��S;L��X���Si�('���%Q����\iq��b��.*��&q+�`��-�4��1wQ'��U��2
�`3��b)&��X���I?:1w�ݩ#�����4,}����������Ӟw�;^���>�;���<M�7�㊾9+���k��(�ȗ�[�m[@33V�p�h�hu?�mlM֎{�ǳ�f}�:�H�쪭H�͡ʅ�G��^L�2_���J�H| z�����YUZ�o���j&R]�=��D�Ǖ?�E�ˈ_��Ə���I�FQ٥;ѥ��BS7*��S�ڏ�m��6��m_��"oBUJˬ�Ժ���P&��t�0���75�I{I��. ��fP�a=YA;۟�d�ſV�S<U,5�i-��
X�B��0*5H�`�*�I�vA(+�2�VT��#�d,-��pWU�ҧh5�B���K6n_'�Fp�������-B��*2����&�,��p�Kܶ�����!%�R
���_��0�s�83[߰3�S�5�؊7���F�)Ed
��#�_��]ό���}�uF�5�w��=�#��w�P�j��/0D��	{�/�ܫOݑ�@�p�p��S�@gjQ��:���!,���7�TdT?A*�$�?)�p� s�s-!Ru�C�f��1U�:K6�����&_�a�B�dN�UCV]�����V��f~�o��t�k`�KU��,����q�h�gA�>�R^������Ƴ�UOs ���2j���+�W9��&��?�L�
���V�]QIE��p�:�b��B��X7v�X�B��m}t�#�
���H�w��DT��<'�����������e�maC'	��i�@����h��9��E���r�Ԧnr�}�ە�;�վf4�xA0��1:�D��)5i2�i�����w')�b[�W2`6~2l�
+���Y$�.������� ����Kl�\b�y��"��/8mښS`:K3��*���_��<���%�W���>v�瓳fun�?!�8O�.TAq&�K(!BW�T4�hzɅlk7�iv�.t��ry�녊2u���h:������:%�q�m��[���R�����X#�����?n"�5�n%;n,J1����0Gāz��ծz���,�eX�W3n��&�FTOQ=�61����`W��B)G����߫�թ�$���Kx�$�p�%��S��{S�7��z�H�{3=�C(�KY�5uk���Y���o����7�������`�/@���[h�y!+x�{!�!`��&�??@:}"�k�K1���@��vqg����8!k4:��e&B��y��K[�pʱ�����a��T{�m�B(�Q�����'��<lͱ?�k���qp�^������{����"�[h�3�1z��u�.J^��J�������ѲS�� �fE<o�5�UN�^j8���}w�c�!�GB6�w�g�1��	���b#?>9�0�FHB�>D�0�o��ꂡP;Y��3�6�^o�d�%��]�T�3C�:b��z{S�P<�#�dv���D0Gq|�W��})[[�[���Ý8���;�>ť�O��f�1�lg�<0}��[���h�B�"�SNq��쥿T��B,}��g*vHFDR���?٥����]��"�,=�
y��b�ڶo�^]^���K?;�G@y�87ij��B"]�^�6�O-�h�orVkE�Hcg�v����\�%����ÒQ��B�s����q�Ћ!_C����i�6���W0�n�M#��W���C4��ئ@5��b�;\tg��C�s7� v=>@�#�[�P�~Չ���k���E�Όbt`���jf�bs�f3",�g��f��f���ģ�Ȓ?#L����Mɧ@V!����?�}����/�7>6�����f�*<�� �?� �pE0��s�v�Q,�0�\���q;�m$@�>��8������k��˻h�/b�P|z���d|����ť5kVŎ�W6�vU��6�r�qD��ɂp5z���.�Š�<G�4Š!SI5���\��oE��#>��<����� �w���Z���\��>�7�4%"_l�L1_���b���U�e �@�����lq0�����خ.�ϼ�L�:W��m��&�!U�3Bm��Y����a@�لԍ5��IX]`CBi�(�������(���\�B$�����G L�:�������F)L>�wW@xH࿞�>y$�U�ਦ	��["�w��n3�UZ�Tx4<{��iNka�N56D�)U�<2�s�G��U��#�T�ݷ]*8�mܨ��Z/ �����8�m~ܘ��jN]B>�����qD(҈�<�T��@�Q58�I
8�7Ͱj���l"ܥ�}b<���_�k�P���ui����6
Y!��l� �3�_*�u�u��O�1�}}��6���/�f��Y��ڈn�Q
?rHo�Y�¤ �-���:�(8+��DJ�����_(NRq$�E�Q�I´V�)^��U�`�������1�A�.�I�UVw*2�����:�3�mL���k39-%n�,�Ū���]-�G�)��f�D�-(r���,�n���,���e���]�nQ���5p�"�m�ی&S�V����I��S(������9_^_����5r.}��a9�c��޿�$�Jش3}���1>F��9:\ ��3e�m���?�bհ�\}�w��XQ+7��P�_`:$���<�!s'<̓�m��Fig��c�'aӉ�H��{��� !	%����#O�Ƴ��y���8"�]�Wj=�1��r͗�Z�#yX�w�(k�A��bW�;��ڽ���A����FY�ܼY�� �ϐ_m~�`���Ӣ��98��k$�P�ק�5��������rN<�TqMTS,,5�~(��������ѷ��*I�r$����c�=�͹�Y,�u#��a���]S��@ﭛ˽��K�^EÍ�䩥_���,Wo�B��=I�x�=y��Ð�wk���	���<ܓ�&R��4��au纘�zл��X_˘-z�F��<*m=p=A ����{%�?�(�R���Tф�B!��*��Z�i�T8bT�|�a�SL���9ϼ��F��>�[�:$W|p�� ��'��#,Ϡ�uY�Sŷ2�{�"UF7�<,$
%Ȏ4���:��$��ϙ�/y�U��[9��/��a���_8���v{߂9�L��]o�t�Zc_wO_@���<I��ǐ}�ԸS�����yÙ�Bf��� ����v�kJ�9$�r*B7]���E��<�Λ��J���jV�zv(�&�����ϰ��D,}�$ĉT��8��)/n*������� 