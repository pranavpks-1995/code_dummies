�M!���!ڨv�����M�dH~ߜ{?��N�<��?����,��N��O�o��=!@���C���t$��ހ
L>ZE m�����7ݟ,W�0�B|�䠂W�6X����`P��A�$���qW�z(^�ҷ��E0��.	G��3��x�kٽ�͕v�
�G���!s��:���n{���05�_j�>���󤒡5W�e�*v���(Sc�������սbD��2��";C��(��)��N�R�bZ��y+��ѭtJ��k�`k�3܀;�Eʔ�n%_�^	�0�=�'CY�*�z��/d�u�4h���qɬ��Aҁ�   � �b-W��Å&){��i�(>�P���1�5���q�0��3������R��ʔF�˒�-�0�P�cPѾmZ�	<�7�@�ۻ�_3��!؟��ͨ`�ab(�)�:���l����,�9���]Un�jG���D����:�Z�L?ǹ�x�ksiъ�i��0�ޢ���eYڨk(����W��bn�t��8>:�.ET�$[�%�d*ʪ{�6 �� �qS�x��L%K�j��..��g>V4ZqC���$ .0�+-����m@����pw����a�517.
!%�/u�_���wĚ�(�ĸ��p���oB��0������Y��|�X�X��Z�]�?�)�W�����~K�E�33k ��P���E;����d#Y�rX�����Eg���f��hthё3���������_�?&�<'�l '��y��!a�a� �(��H�^��&U���E[���������!���"�"X�F���*��6�Y��F�L�p��|��S΍*�!TD�����#��  W#��w����F���#S�c��p�G+�V�XX�Ä�^|$���5��N�2|4ݳ�:�8έ���c� �9�L��mx}��H`�PPyM8�A�H�f?5}�r3e\R@    !���FGH!����X� h����~�����?���^���t;}%ؤ�����'�y����XH�'V%�^��ww�7M���N��
�]���/��ק=~�Y�^p��U�=|'��-�q()����GDw�-Q)�\��>`Ec���HB�<��0i�!���"0�bV= ��	Y*Tj�����0�rm�ّS4�U��}ʙ�� #�B,��`EgG�`���{�$���f߯���,�c%Z,�9et�IU���Iy����`s�
˳� ������_��Zd���m<�#h