�U�/��5�宣�쇞dm�YR2��/��������+����T���w�����viDqb����V����BH@�`S��E��P���|�S�CiA봏E��W����/��<o��xU3l���Xn��
lH)
�����`�9��7�by}�h��Hު�6�x?8�O!D�Pd;)Q[77�׷DS2*V���W�;�&hım4n�,�ڞ҄^9 ��������7
(�ja�VlݹQ!={��X�?ӽ���{v��R����qz����Օ�+�%�B�����ΰ4�@��v]����9�"�ՙ���n���VmS�4���&O�	~ƤH� �b�M����1��ҧ���o�JX��i�ñ�Ʒw ��-��_4C�s��u��w�c�V�����i��Z,`_�8T����?���E��_���'0��1Y�[G����&�#�R�t�Y;��'���<A� n�Z#�.kP¥����v,O�ר���ƣj��4?T�~ǳ�-�32�O/Ъd�_�^�f�64_j��9�����J�=a}�$�>��z����X�,�Q�z�k�P>�M�(*3���t�/���1����,+)�F���Z�{��Wjj�|E�e