g�Yx�|4D�y�����F�YF�p�S<�uA1�"��[ǐ�$'L�v�%�2�"E�٫� !%E���+7�Cqg!m���*�t���~�Q�$\��᧽�z�`�	�G	G՘i�mқO��d�HM�������У]D�º�_�"J@���{�?s7�F �B: b��E�#b���:0���_��V�c�CAIG��} �!�,�Gzv����v;<	ynU�J��f�AS�V��sun~J����`��[�wMQ����:��0:�]�B"�\ut�������1S�Q�2}ț*�����6���\��bIf�k�!Oho̼��Ѭ77�@{pa��ˡ~r�-�b��6E��� 9*��@@��B4�J�͌G������M\J�`&f�N>�+X�:�y�"z� ��@��;T%$�sĪ��
���!�g���&�1��z�Ա�5:�����T�k�Cu�O��2f����^�Z�f�>wL������/qy�������ڻ�̍��C֜�]+E3��L�h^̪������� �eA��ì���iN�?F���.���q K9�7=�W~�M�xˤ��ތ�H��d95�)�~;��P'���D��8N��i�r�$��~A�C�u"��Hޣ ^
�  �  ^*��]!\D`�zs�y`�����wU]��N�f��
�s_�"v揇�8����@"�����_V�3�8�-���g�+0C�N. t��$������G���e9:�KQ������?�Lu#�aB��@U�bv('��<�~k�_��x��u��Nڹ�HE���������V�C������=���P�UL���u�$��`���7��0�a4աHR�PT��l�HFeן�J�K��Q��⡸�]~z���E�ۯ#�T'|�P�w�t�P�,����{���+M�� ��f�+�{�Of\NX̵+2���͠x��� ІT2SѮ��e�������L���K
��XG$�,&��G�|#t5���:,�ŧ]�H���~�M��לUv�&0��K�%��.��?�F?�J�?{�8r2�y�&�0�_���̌z�V~�=l N��6�Ǥ�w��z?��!�>���x|"��@6kg�D\�Bƫ(fP�V>_Ο�x`rZ1�'��ky�Y����$�_�^H�:Oe��  nOE|r�?��S~�h��
�3l�����`���V����u����kқ����LMMQ�v���(+@�S8�X���
�2J{�C�j�B
�\��2kR�s�S%�m�����>m�K�_�Ԭ��GW��������:���R�1V���(���K�yظ���Ō(?֎���J��^��ES��1jyx���RW������Mjy����ȡ��SY �ID'��L����� &�q��Pv��.�B��P�]Y��T��r�.�%��M�hGj%���Uz�3wM�y�r�
��1	x��n�
D��,�cPK����J��$�DpCO���*%� 9NxҶ�����f!O���S;!܍�z�f|N��y-���,˙��r�ees�l^�hi����7B\Az[��X�i���j�_�cYa�Ͻ��*�QXN+���l�
$��M�bT!����X<�U��M?�]�_08e�Pf@CT!��s9����łm��s���W ��1ϴ��]i�U���Fz/$��>