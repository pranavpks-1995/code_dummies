�����5�`�0��f�̾̔��|<ܮ��a���8J�R��V��7��g�k`�l�;�c}�1�K�0֋�?�XT���r�֏*���B���?tK�]�.�)��Y��d;D��L]�/^$VoĠ�գ�� '<��M�p�R����]�g^ܠ����3'.�u���t�|��@��VX�J_@U=�g�A%��**�{�bh6έ�M�D؁'   � �F�u�!j�O��u,l���Or�A6��|G^�ǯ��
��+����e�S'���1���%k��P͗��<I5�^���AY��N��xo��$�?֡ڔڭ���o��B ���9��	�� �t�h�jU��T[oˢ��n�E�
!��u�fj��=��v����!�M!��,��H@�1!fA$ }:x}::��@d��&
��<tM�����HJ7Ht@��𞪟0�@(�|��I{�Yz�w#ccm<MB
u��]Y�<��\b�/I��l�oCt�m3yQH~�&�u�b9S�)��B�ζ�6�E�E
��ء�[�@4��]�4�2�CIeU�Hv�B��s#�	��l��^[�������4D�5�FC��}�#]��iv:N*;?�&��!�Pe��O%�`R��� 9��QJ�����|\M�n�m/4T�������C�ŞH�E��4����6q��.pJ�Ǒ*A$���ķr�m�TF����6`�^�q-O"�-(м.J~a��D�ﴐ��EF���o�z��s�uY�:��Աzjus_ �MZ��dH*,UZ�	���=���YS*<�`������ .Q >'�x�5�Ҋ!,�2�h�

,@E�8m`��Ĩ�L�`�US�R���7D���s��_��hoq
���E�C�O&~���"+ǧ�D��_9��k��gH65>��H�,�/<Z�]շ������\&v�cΨ	�B��U�<�`Atw�k.-���	��ҧ�=`]�?�D�h����I>����n$ j��Qj�',]�	�[z��W4�=����j�B��̈�=�*����֓���%��}�T��߭��Rl�+b��N�O��	UP��{^�	��`~�Z�I1�,:0S(h0Ʈ7{�Y�` (;[�v`h��fT�Jb,h�O:�L$���Ҋ��+��<�iNAv֩�{�҈E������V�n�b��D-|��@?���w�=!܂lV����k�xR�*6
ó]{���̿�Gܛ�2�_�L�{ ؂����X�V��Es߷Z�ԇS�f��#UL �@���uQ��7�LNGP({Z�S��qo�|�Љ`ݢ"���I"Ѧ_�%l~͘+n��@���~uT��k[,��/�Q�Y�0����L������vTfMf:�o���q��-�IJ�N�����Xc��7羧9,��$�?g�G����-��d��o��b_���B��z   � �-���ún����٤,n徶$k�_Ğ+�T#��l��$�_����@�+����F�\  H[�@L�/�T����.%` �1��s]A���=�B����As�~7m��a�ۃM���d�AFe`K��/�Ѐ���T�Or(6�;�r~Z:F�|T�b"�K�� y�v9OH�0��o
�F&ux�� �5����g�јO�?�cV�_����#��t�u����R�f������:�����ϥ���_u�;P�Spu|J܄�}���`������)����]�B�����n	Muq��e?<BҌ ���zJc�K��M��R��\;�2ɱ[RN�����r�Z8�Z��WL��Z�xIw�k�����?����o���L6��B��8u���1\!(y��$.�����+����p�Ů�< �EV;��g+Rݤw�6d?ڎ�V?V�Vz}7�u5х�4�~���H9�@�G+!'%00�&��X�Y����#��Բu(vgo�]��v3ik�O��[J����,���y�9gu�,�\u���YsW6�S2�"������i���z��Ij����Pf�I�Ն�e��N���{�=��w���PmM�G?|��@݅�4�~�a"n���oɨD'��+��Z��<��E��	��������!��A*!M��V�
��%	�d�n�%^�+PF&�Ɉ�ZX͒LT��1e������սښ���n��)Ô�s��k��]lX振�b��-�=��V�#���gw��GW�?\-�T�qq�����跫+�I���$�r�� A8 ���~oT]?w7��N+C׺m�B���j��   !��8������� 2�G�F�=��3�r̅g	ݖ'�S�,���	{h>�P��ON�-?]��su4�xP���5r��7{���������'8g��ZtQ޹.g�r��nvWQу�X� aS1Q��2�ɫ�	&`�! @X R��8M��!iT3w݉, K�i�a�
�Evi
�^�-� p!��1"�" D@ W	�C,"0,nS�4ٙĶ��+y��	Kx�~�ߙG��r���j��.󫵖���D�XgM=��]W��	ůRd?��PCDY�5�F��g�B@�m�j5���[R~��3O�7�Ɋ0[�!�����f
 � ` C@9���Viݪ���k�؊k!Js�n o�5UK�S��l     �!��0I:ĩ4�)�)���� �\l��t�4�e��;5�"�����i�������-��t����H��0Xa��f�cq�@��uu�#W��匿�7�^|7���)\~]G|����>�yR��T�  H��h �� ��}Gga�P���4����~�*I6��   �!��9X�" �B  24E9V�ߨ�`"MŉP D"�N5��*ӅL�Y�R�Ql���"D��U��O�tD~�����87 �7\7*Q�UNa	���h���{Y^$;��2D�)�K����R`$�d�`4 ` Yua�9u��WF	l�%"JTŪ�	�f�hsw
d�j�0    �!��!X�`�Hb�`@!��-9yh�ib����=W�V��B/�EU�8MD�1?*LO(|�\�,}��|� �#À����0BP���ӯ�����2�������'4v�Lؤ�:���K,��