��)�n�a3X�W� �������ߵ�;�����II� g�]�#��U��Y-�
��w�	�0r/�G�> ��?u����<�45 h�o�CG���Kp^�ś]����q�
l�밞ܸ�� -�ݚK&*�׃ϙ2�2bĀ�Dgdk��6s��2��C����8p�@:��4�{���8 :�}�i���_�S���ʕ~R��A�������b��G��غ��顙m{+�~�&�I�r�}���9c�ݬ�-7�C��!�f�7�lB����ػF�ќgW�N��ĉ-�yɏA������3�v/ne<��Ү_�g(L�{��Aԧg��
#K�p�k�h�bw��}<N��ڧ��`pPX{&L'��`��K���k9r)
��ͦ�j ͧ���ę������J�P�dr2�F!����;Ǹ���]��+�[��^��������n4�F��&������Z
(�B3��d��U��8�i��N1�I�)�L�	�k Hxp�wȌ�fA5Q�����^FKbԷ+MN�m[��/V#�n���s�|�3�^*H��`Xy�.�E��fc�jHs�h ��3��f#����y���҃��M'��B�S���σ.D�F'�Z���/����tx���-Woyc^{(�ϳ��X�_J�j����\��&N��v'�\M6wW�]W~��Ơ�`���p�3A��I�1�~6j#z�{�.���#�߿M}o������31Y$������֐Drd^%�� [d0�'����"�����}�M�;�<:v�|53��h	�3A+ȓ�Ք���"��"���:둭�&=!B]T%�����ڴN2�V�#��d�'�7��ƳB7��������; �]]#�[���n^�ti��6��{41��Ρ�SƙT���Y֞=�5j&'�����Yw��O�� Q���-O�1�s����{"M��i��,m��	YX��"��ǲ�1�P��w�e뾕Ǽ[�Ƨ����X�O���j�;d�HA'i���ן�
,Xm�4AO�Χ���0A�+ZaK� ��6`�����v(��W�;�R�b�zF�E��VG0�U{��x�7��fF���O���m�?�uK�k`��g;�d�n�K��Gne�=g�d� �vwt�A�d��ơ����!���ci��Bٕ�3��*��l��7���p�,[ ��m�`l�SNJ�0�3��KZ^?���E4 ��ᕭxNs����e=�y�QT^+=6"̠։ ��. �7�� �#��r�v #~<�+Z��N�ő.���Q��ˏ'