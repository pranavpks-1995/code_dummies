����Ǒ{�mL����D���q�f���[�kX����%�AA���|���X�j�/�Bw�?��$�j���vb���EK�˂�������!��=f"��`    ��]��?�=�k^�9���W�`� ���`z<��7��IJ ��V��%.�t0�c2n���)m��rl��i_似?����{�R����`  6 *G�*@��쵬��*,��D08����ǟ�����9@ �.��.@zB��)
�(0  !��1
5  
ΊV _���\H���e��@ |���S�yn#W�`"�2m����j	�J��`��i�X�M�^���ʖ�X,�8�@�x(��.  ����V��}�����V�8��*?ib$[t����7�/е����& ֪�` ��o��T����� h �!��8�/AC��%� �.�%b���e0e���nMr���أmi�1������'�P��a쇎w�,�aVHL�-,�(P�r+���	�40�5��kX��4�Ao�q�&��@*)���r6�,j�RȽ\�+:C�iR��B��@p0� !����"� �� �`5{4 �`;�LZ����R|ae��`�����f>��4[`�QA}��Y] �J��%�kD�+��"��H]8�@���	H�h� `,h�l���d}�i�����v��.�_X����zvN�&dp4�U"�F��  8!��\�&K�*���� R�q�U�b�J�߷g�{޸9Ѡ��)V� �ԁ]$d���InK������TX���W�	�X�Q3�ӡ��9�`#�R5�"2�D�x!x����na�s�@� "�, Xpfs�M��o�����)]Z	��ʆ�!UH�c�D�  !���E���50�f���e���h,�7��@8Px�A羓3�.K'Y3���������Q�8\�"�P���u�R����j^�<�]�+�~�9R��X,D'v��!(��� @w�r��)b=j��mh���!s���1N�gl�^w�%��H@8��^����0 0!)��5V.  XE.������H�"k�afnU�E�Xv̰��*�&�FQ��Qj�
xm���Z���n��6h�ZкB�����0�WNtYC���}��&�N�� @Lڵr`�1�X���ip&�9��a�!_��3���Wp'^���"Ƃ�  !K�H1>؏uS^hD�/3Z��T  V��h=�|{���J^���X���7��+��4�^�G�;R�ȨQ{E3H�'�I�-oh���=�׾����Zh e�8����~~H|�vo��W;���D<D4$ �<t������[GSkݽ����TD,�e�L�a;�C:&�!uID��J  �E��   �׈����C��<M��ƥt�V� ��81�
?�P�%%�c��*	�E@rk.|V�3�2�.�O�?tg�A�_�S��?��g�˨�X\�Cd�{�Ҁ��m�)�}�T��{BFx����n'9[�~	�������$����W;�S�r�#��؟-�Ŀ	�1'����g'�bd�jo���u��°6��X��6�M�	M'n!��YEf�O��g'����d��@�1�RqG'$�%<V���b�d���ģ-����r�c���ϙ��G�:z��[#u2�u"|ߒ���8�r�i �R�-`���8Ѽ"�M#���ݼR+���z�qX<���vb��A�]�J�Q�e����n���A@�]H��Y���0*<���g�c�>��`��║"�O�B�(� "ڳÜ�K�~8���q���T��ƕN�徃4�
w����^)��~������cJ��ϰ���XA`������ʒ���U�[Ð(�������
깦���~��_8D�3��/�ೃ
�+I�D��r9�+t����,�}W��t�Q���:��V���(�`��x|ڍto�d�>�	.�ق�KU{�;��>��D�ү'0�P1֢I�@�;����M@
�O#��䠢� �p8��w�uZi��cfPC;�#Ҷ|�NuM��O�4#B���d�@.����<kcL���!�ڤ���0�<�$���U�=�$��x���C�fA�O�Ow^�}5�zC�*�9a��[Q>DM�%�|�ժ�
r;myqI��$蛵�K�pΟ.�V^�eL�l9�'���Tm���"�k�A�qk�!���5�{YiN��Rֻ��G����Q\�n
����(wO/@_�x�ۡ�9�/�O����J�#�YIM��}mw�'�Q��,���3Jx��_ֻZ��OԬ�is۸2�?�Y&�ؾުI�3�h�k��ڊ��h��