�5������|�������5N�c�?)���S5I[��`��귅�k�����f���j�W��%s��p�N�v�Yg!r��ׯ�,�3��Q�e�,��C3��c�����4��&�@ҷ��c勨x����9cȶ�R�>�p�	�$�/�Ng�ΕI�����v��ؕX=W���m��C^]@����P����)^��%c���TLT��Wg`�IpB�W�è�g���hn�Y8"�Q������q=�@U[w�������e���H�֦W˽�G�qZ�\)
۪��1J��sX�q�K\�&���M�z�V�]���̀` @�.�&e�HM�&n�r�~�O$��8`Q�z���_��:O���%�4h�+���Y��lX��s̽�s��:�{1���Q �n���1w/�V�����ߨA�J�P��v!w����g<��7 �f�DXwH�������
*��	���.��*$=�4l��ȋ�n���Va����Gi�m
�P���)�	��L�<���5�H�:�������.(�BJ��C�4�T|W����U�;�x�-Z�ˡf6�	�ɲ{y�{j�a^��/���ԯy�F\���B�>D{�d?�B��j �O2�@Uf�3'����9����m���p�����Eڠٿ���:W�r>V6k�p�'I�B�ĞF�Dd�J��g��cJĊb9Y�6/2���}.��r�=�!{
'����%�L(�Cn3��X�H����P
�pm�@S�ډ�������/E�Q�@K�~'udq_q�j�[2ԣ��4hܮ����_~3\�W�ؠx\}�x�g���E.�)���_P�S�f�ZB��u�rY�ߝo��lY�E;�e�C8�M��/alD)�f�VS; �p��n�+�� ��a��gq�@f!�;n>:���U�^=Gfm����������e�.����<��/�d��.����t�p���wi��2rn6ի������y�q���ϭJf�:��&h�T��da��]A�H��ZY�"΋Q��5�\�68��6�፯�7�
���K!�Ǻ)%�ȃ�f�ܡ��SQ��Xr�����rCH��㌏{��-W��E�]O-�JUX��Θ�[7Ũ��b��\��c0�&q���=4^�� �Yr�1�!�R����ա8߾u���D�/}�P�x��NG <��MuH) ���r	��}�x���?��VS�j�ڸ��/fȁhb���"71�F��q��ѹ� O���cB������(�;5����L|��MQ5�P\�eɰ�^�CC�%�5q�)<�J��=�8��,J\H,��@X&�`�
���ؐ���w���?L0O��Bv�/�:������3��6,�5=�.� ���k��#�?�\M�I����]^�������/�������!�sw:�5���A�`� �}1�O��1׹�V	r�	V�{ڿ���L���i~��\�B�s��p5u����Y;���Z�!_�V��(>]Ư���&�ohV�JQsSC�>�~G����_1:l��l>�@U��B�>��b��s='+[b�?��/��'e�������uI�	dlX��} � �4���(�'�@FN3�x���Z��뢿�5�·[l�M8z= �>�t�¶�Z���C���q�uȍ�l(�4�Y��5H�� o��*B�ţ�)��R���Ds�"��W��ML�I�5��$�h��p���p�Տm�%�6���Of&쭓����Tݗ����%�'P��3�b��B۬�Kї�ɁϠf��������O�>X� F�z+����;=��c)��T_N μ�mH'�A�4��)�Ĥ��*@u3$��v�2���,Psn����c���_XT�猢пRl��5�-i��抂9L\]#gyZ?�x�����q|��d��X��Cן�e�F|�r���X0"�VNc�-�5�cz�C&o튜�Q�ꈻFs�!����cJx�,����u���@��$ֱ��/��L3���h4�(��\X��"XZ�)љ�+��8q*�h&{}��E��-\������jث�4Ur|����홌�,b�'@�,R�T�Ř�hᆾ*MS;%�3_�����몝��4�4J�͚��8���n e,�6MG�R��WM�m����DJ��>G���^QG	cc���]U���n3w<��*�1��½c��#'��@)Jn~/(�1����x��[:�t|����LI(�Lqn{�'�F��~�������J9���X� �V�;�`�����p�r�