�i�\Z������M�66/�?�e� �4%	��z�B��jWV��S�h��ڐ��S���ql`k�X��l�X	� ��ؔ&��c5�p�ͧ�� �*~�h}O��~؀x�ɮt��F�k�LT�<	3�&/R��ڎW���B��0�S�M@L&d������ŋ�(q�%�"��!i���;�X��xu�уV�X�oq�O@ͪ��
 ����ݣs��	�����)9,��Q�X\6Pg����w��.n�r��y6���"�����z���z#4|V���oc�{�ʒ��1Z�0(P'L����LG��Qe� *�-B繗��g=g��3l9��i�Cݼ�Y�.�0l@��ْ k���:��S.�<����ʪ	5bdk�h���VE�1Wr�(���L�����Y�X�!�9=謵Jfbe�6��?��M����=� 6�잺!�ol�W��2�
ߑ�oh�2�UBb��5��:�N2�1�3S����x�٘#��y�IV�~�a��Y.S�l�l��\��ۑh�(E�F̴�}=��5���@�R��"�@��`�?1�3�uDj	CX2��:�ORb�ܕȋ�i�������Y���y����X<���,.������]K�V������I�-�w��N�h�^-����W_#�GΞUH��;��X���$hl�w*r._�����G�G��Λ�TB>n1��g��vv�v�#u{�O��Ƙ�-ݞ(&�v	y�R��b�v�^������庲m�dD�B[L�n��ps>f���ɑ{4��S��t�@r�~���OL���H�����V��@�[*������Cr���IkO���Bo�!lkh�E]n̓v�~�om�\M�'"���u)�V���jVQ�3xRL�����,zV�r���3Ztѣl���v��̽������)�&5��ǩf�z�K�v/� �x�)=���T�ӓF��.l\r^���(3��V��-U����i�j����9��#n�8����s�����v��㰫s{jŊ[��Q�GA�*�mO�d� 
tK��̶M>A˿Czy�(r��E��/�ѓ�$��]@Aƨb���/U̔l
�9�"����F�b���)ؙ�P��
[-��N��Ʈ�s4��(�1�<sb�cP���=�AX*zG��N:��;��|�b*^�)������/$o����N_~�BU�i���<��w(���o�����A��
  ���'RW�c�`���'�.8p��Zy��j��X��b�E�{�AH~UoZ⇱G�" �Y��c����GS�51׀�y��;�(�,E�Q�JQp�V���q=��]�c��m}N�ǵ�i�[ ���#Z8����D-+غ
�J��G�q1�H̪W� Ae��X?�r��~ O���S	}>���Й���/���
,� ǬZ�Z�n�O��r��v᳉�H]��#�{l���\�_�?��a1{ݟ��a�<Ί�/���,=Zx�G\�W2F�T]��t�~+d)��8`����g���~!�l_|�;�s�$���ڀ�PFw�Ȫ�\�UE�tBʹ���y!�Oq�Ƹ���-}D��́&i�E�/�qlʥ� ��i&#`W��^�Ti�-���Ș��A �	�   � ��U�c�}dcL�J�KA�N��M��#,�H�ɂ�����@��ѽ͍Ӫ�Pm��৶}?�9Ow�0ݴ�~jٷ[��GKR�Ҍ���L�}��«=���e�
`B-� 1�_p�r�8�.7Mk_L��Si~��⊊>��C���J��/���-�ݱua�4Θ����/�vU���yP�d�m<?a��l��dH�_0���F�mm=-�9�hny�<��Xi�n���]�.Kuf�hzZ.l�A�	�    ��u�e�Q3�eT�*�� NhG�w�M!��y'��\p�15Y��{J���y���7O4�4�����D}�/��#�9U}n�ݛ��O��2�n�B�h6�9,�){�X�f���S?p�.�W�.襝�ҟ^��\��Ψ����>=�lu"��sz�{M�U�+�ä��VN�CZ��0��z;W�~j���$	���*
҃Y����~����I��{�w��r�͎�'����~0�p�{\SS��J���O��A�
D    � ��-����bHek9P�8Յ=���H�H��3F�0#O�>*�2�u�lNy�]J���eY��o�����w�^���cb�TbF�M�M�H�@n�"�ٙ�>��Y���e�H�ʸ���]��}�;}"���ʱ����\3�(.@t���VB7�Z�[��BE��HPKH�?� PuW�!����)+r�m/��o@��9�"�:�p��u��J$вG�bNJ�Q���@��k�c���/s���D��
���������!��A���((�$(�d��!�@���!9I��F���6܇[�v��Z�_߯�'�UON�����(���d�塯ԩ�/�O���㗘��N�(K�ΰ7ƚ�]�r�������q��P�>EP�Я�H��E\-~����    !����!� h.��
��xT�F�p*�SF���BG�>5Ɯ�!�߾c���O�P��t@���u޶W���V+SCJru� a�@k�hԂz{n�n��f��f�̻+Я&�V曍�:,�"4�C��m%�B`
 ;L����HBS׹gg%@` !������$��"
R��aR���ϫ�"�3�\�������G�kVD��5����FW�@"��@5��`��0��r�9 � e�X�WW�֦�]7�z��Ǆ�N}`�`&ȡ����u�4��3ɲ�a  8!���-�L��� �L�X"�;��ҁ�0/W�T�`�[0Z��}ohB�Jc�.5���/�|���������H�y}05{���D���/N�y�}VX���߾q��9��G�7��3� ��5'�a�%���{� B��p�����C@`!�붂hr@��0<Z�U�V���;1Uvp0q� ��|�6�@��)���u�r}oF�k}���ݠ����[�)�l�+S�,�M�)�g]�ˡ�o����?�1
|X�Y�檒=�$�W��$�����3WQn0���ǒ�bP��A]E�i
�P?o96�0   p!����ݘU�e,'C�'�
���|�/W��G��j鄡�i��������0��������5D�{�o��t�Z$�fU�HS�o���s�̀;�ֳ>��_q
q_��m���D��J�*&���0� M�o[t��5y��-   8!�����S��T#02Ֆ�� �.R�w��"�?q�Ӹ
���Z�p0�W+��s@\�a���K+��_�{�L�0j�;�E�����y8fk|o�����Wf u�&�f�?���R�~�����Fs����9�gP1� �5  ����	m����	��`  �!�	�Ȣ��Ռ"	vrpa�Ǝ��2�K�����綐0y!�>Q���ii�Ԉmc��T�f�)G3J }�Î *��D���HK�9���Y?��荂�F� _W�~Vr�z��gs%,����`������ L�C� ���W�H_����}���  �H��>   �Ԩ����C�����܌�S�T�0 �H�`��o�u_����΅U[����᫁*���5�
l��X 8&Nw���\��bq�;NaM$l�_R.�싟�h���teyܵm�i�wְ�T>�ہ�M7T!uԾVC�ߗt�$�%�b`KQ�����};3K��)��$l�X���� 
9[�x��9��Ǣ��;f�-]�g�Mc��Jڛ�6�����fZ"о�u�J���.	5��栦��;���uN~�m��v~ӗ���B�1��_��:H���/�dө��zFQr_�,�5�8��k�r?�z��7+�(�O+��)Nj�߱4�, ��{�ة��D��Q����\*�8H���ARĩ0Hq������~.TQa��ջ�	5$�z���p6�j�yzϼV5�l1���S�� rB?�x�S]�6�~�b�6t�xm''��1�Ɩ��B����h�X�ēD�r&��2<'�������1� H�9��{�)�=f�IJ�:��+5uА[9����U��I�y�������E�u�X,ǂ�_�@N�	��"��[�j�cÒ_��ol�$��O��+Kl�����0̉�A>A���m4F���Z7�s6Gz
�k��6C��z�W��"�����f�L��ڰ9!<8���LT�3c�Y�FM��lfd*<r��>3��cV�'V��C�T�x��`J�䃼�G����p@�R�HЉj7��{��8�]�0k!uC�!8���ʻ\��[�^>�-�C Y߶�Ѣ��K�|�������P�i��m%zMԻe��U��.K�Xo�/2��q��� �@�"���M5��/�'Pۖ�i�������=�����������Kc���:�?�*E���P�!����
 j��/_��*�ì}L�?{�hю�i�)Ga�M�Ҏ��㐞[>BfD��n,�(6�6=բ��#�<�La�	�l��|�������N�P��@8�r��l����o�R��M�hm=>��Ѵ�M�L�H��)�Ⱦ�}y��4��Rw-6vIR,'��`�v�xg�rY���jî�4�J@|��J�G��.wd�`qX�*�q��=�$��RV�s���%.`�.��QxN�iM�.�����1r�C�Y���w�1T�$-�� lg�������� ꔗ@���g	��:���+$�,���r�εc0��
�J�nK1�Lg��?	��c��f����P�
�}�	��d��|[K����Z�[Z �.��P�c~݉���Z�q�+�F����?��yt�K�y��s�3>O�ڪ�1X��Ш9x��L]+X4�#L��]t�I�z�[A�jGe$�iq�ȱ��V� (˸�`r����j�MA� ��3�Q&h�zШ�89� �_c�y[J�\��,��6@|������'�O����yx��} ��X���z���#�(�?�1��"Ց�^�o͚���oL�7��!{n�O'�����������Gk�+����(=����`�D��HZ�U��m�=�S�p3V��ʂ��J���1Ʌ�m��L��(���k�	mKI�ex�ǒ4��b�	lE4#��C�Н��X�{�ln����K�#�rx\���w�(]�i`��Γ7��S���A?���� ���	ɭ�CG7�yAy�ڦ�a�$|��\�`D�w�\���dkE�.Id^��#-S\`��N?�^��T��^]0�/o��!�HC$���vm�2�����l�]������  #� / MėO���Bj9�%uؿ
gЋ����Zhb�؁���;�ł���l$e�N�O�K�?���{Rv���%(���wE���Ɂ`��ҩ�ٷݙ{�l��c��Dg�u��͉�_�Q�w�ŷ ^���ٕ�-�F	��t�2�P~�p׃QO�[�@���S[�O� /�t(f������w�3u�63�:�C�ϼ��.�{�����<,��:R( <T����ț��"��6]iU�| �?wk��B&@\o��
+�)R�=e�̺j.��8sta�����S�ax�k�ml��?oN�-JE쓬��!>��^�=�>	mߺ_� �Q/U�[jU��{��j�T�Y���\쩝��}ߖ�n;(@N�s����6gŭ+R$����ً��z�m���*�$~��P�޹E䓅"�I&����[��c%?[��y��v�q��R����4ԣBZ�
�  R�b'R��c�vd�j�4l����ܞ7�iF���E��ea�㿂j��=�deW��)����j�K	K��@��m��3C��4��u7٭{07�������mRo0
}��X\�9j7S$��}�����B��,��MEؐ�pt����
��T���;�!�r���"y�%5��F�2��eY�/1�g���gD�ؓ����/��`�� �E<�P��9C>5�@pǟ=���f�J��V+z]�����f��B��8EC��4���[S3�4(��ȭQ���"�t��N�q�kc�=Y1��̢��3x��5�ŻKq�=���P��?߸u�X������*��AY.i����ϻC.�4�æǍ/r��jKi�!