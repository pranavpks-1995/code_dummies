^{Cq0��an��������e��E���>�w )<q>6���l�6�4�>V@�j��T�B�sӥi�T�_�ӡ��4xj����(�.'`H��X7�L,Q�)���CB�`�m�>
[v-գ�+�2c,�Ǩ�Vɾ�&��d��'N4Q.q�g3x�CP��T�����U8@�vډ�Ľ��@�͒��Tm�������|x��0Pt�Ng(7lrp�� ~��dk�fCrw@����cvwC+���p��* f^����	*֕��{k�J�DH��u�!o��5��
����38�Tn9-մ���
���و��'�|G2�B�۱����Ju��R%W�(l|�M���������ZL��E]�Jͮw�©�9-KH����2�
�n�'�O�犽����ϓ�(�*)�u��h���(��M?���N	������$�wM�v/���k�\b��5�Xb0L��.��Q�����W�݈���Jo�G{�C�D:q�w��d����t�d�����z�9����/H����2Y�m����<bC���m��[� �9��lu��t����\��u���G���W+b�e~���u�1E��n���V$�H���U�GꆹǶ�#c��OO׈7�j�lz�=�x-#�/���_W��wq�m �O�Br����8N)�������f:$�hY�u^��jE��d�w��mr����T�]eR����f��2��wKs�P�!�x�_�7S 1}1QZOT3[_`ƪ���_~a)��	�sg��\���?Lϼ>�����������������������W܃p�]q��v�;���%�3��u�f��-н�;Rqʒ���p(i���C�i:0��'d<����GyP�l\d��@�w[w(�wc���&���)M��4F��$4c2ӊ3�Ae�����H��B�㱐jv���9?�oz֯°%Vaecv���z��ګ���3������3��1��I�YY�ZÊ��ty����.�X����b�dUK�A�]y9��h����m��|�4ˊ���aXK>j1��	�Ͻ�'ߒ�aIR�l���Aހ(p��f����g��90 G��UG)Qn���3���x�L!���:��G�Gc��H]jM�|6M��E0���F�h,��}P�f�W�A�,���Bs���g,
�5�%)�E��PD�:��O����q�� :���.^��i�3�Ui����mg1g���n�g�^�E3�iHH̔�CH��>Y=}@#�NI�Ͱ;��;2~�ҁ�U���9j�i��T9F�H ��@�Iן�6,�����ϝw�!e�� h�B��G J�_�?yN%=���y�d�״��-�d{h(�,ZΒ`�Y�*��
ME{�;�f����<$��^X�r�p�Z���dB��9P�:��ܦ��V��R'#*�㬐�a��5˥�T���`��"��G�lpˏX���`\N�@[�'h� �C�a
}�B�`Y��Q��0��v��@� ��PY�Cl ��myuK�<� U�S3u�sBa���� �J��A����D�cff�p�*�����b<�[���N��7b�ܪ�Ӧ����0�]�u[19D�℠|	^�4�-�4�&b��aF���Io*���K���(�,+t�t_�+<KA��5��<�LThӪ��#_(��y�/I�õ�d&�x���D���l3ciG�ZL:����W+�AR���-�hL%�3�^��0�^�S`&��0��Wh,�T�O��F�ԑ��'�O}6�.d-���&�w<²�5$��E�m��֫���A0*4+lM�k"�Z�{�\�x������P��dFt҈��1A_;�;D-^,�[d7��'��D������)��2�M�`b $R������e��Ux庴H����E/�fO�`jO��<��u�� �-��8> ���m�d)Ƿ���]o��8����K�i��,�K�μ9r�d䥉�m^T'��h�#��E"�6(�c�x��i~��g5iU�M�.�%4 ^<��Dv2~x�}�ň����ڸ��Nԕ���w�����I��0�A�\U�+�u�\]������R�`]�t�b���k�=x��~�x����ɃL�k3(�wV%H���qE@�3��v��F�⻊��p-R�q�'����8��/��sM1�d�]����+*:i�k�aC�c�L��?D�M(\�����9��4F�0x�pJED[���?D�D��f��{F� c�INj"]��y��@����Y���5�6pE
 �NA���s8=E�Z �9/�@h����`�#O~aƩ��\���uX���uH�W�xh
��DFaG�ճ��@,O�-ek������?Z�6���9��kkN��"�4���ޡF{ĩO���ك�#
��&�+�X{f��Z;
� �_F|�`)F���p��cQ�Ğ�xxS8����i�y���!6f<�#�)��1�/p黛��݆2j�i�+����|Mԫ�a��Tm!�#�=A@�rq��Xm��	�O3� I�2�8�]��9lei���f��L�b��as/���{v�lg�b�S��X%�D._`����'i�3���(E#.�\���*�Xj�b9js�6 
�c8�1m:"-��$Y�hٵ�$c-y�R9
b!��A<n��L 9G��fz�|�pאu�ŵsb%�o#a����v-�C�s1qC�']㈌S��90�AĤ
eB��W	8o�+���P��@�Q�v.ٜܶN�d���:�FL� �T�D��B����懹��1z���E�*)T��6C����{�2���7�-���erH怔O���Vy��ߦ9�0� Rk��6�@h�T����փTՠ�{e��������}tQi�����i|j�<XUXQ�߸?(�ri��]��m��g,h���}=@����M5�?Q�����i@i��7P��C�.an�#!�P�*����x=��0׬x)x6W�b>d��v8�+B��<�;{K�	��͘$$E�bW&��ZU�t,^۾30�^J��{���Ȳս0D�~Z�e�>�>���7M��K�a�������(��
GO'j�̕��3b��/�.	Fzc���V��������`
������]iR?�-�]3hG:}��u�