K�K��w�Ӧm�T�]9A�#�C�%Z� ����A���>s�»	��/��~;��X�B�F�Gm�4��S�:cf��Z��+z4Q��	��g���Nzݐ��DP&��W<�?�x�rl�6�5�_�\ײ� \�L9����P�=B�t�F[w:
��6�`��<�)�;De*�L�A�ƶ~צ��b��K݉x��q>����D ��YQ�Ń��3�P�����b5ܫdG��� 1���`:l�g���
a1��.�6Bgb���v�ބ�6���m>���#���Z��cl���axt�I.ȑV���A񽸿O� �a�O��5�����MrU�.�tH0M@�d�k�:�1��E-����ی1�M��'���|2ǅ;�ȴ��2�J�=JP�`�a�y~�����m*�)��J�.t�hT���̀�2��'���`0.�u��� �S�⿔�V��i��*��K&o
�)4&(g��!�a�E]A�G,xJ�^@�gl3"���m퍢l�H����;m�ؠ�`���	Y����dF�afqWf���gW�\?]J����WD��R &,����!�"����{��~�$��,|��*���d#&���T�{��B�x�������O����Z�d��6��	���I�k<V� ��BT6�v��J�+g���ү��2@�����gw[�HW']��GC�uK���H��>�Db�f�aZJ� ����k
��߄@S ��O��x�O��AQ*�˸͞�?�)�\�b�n�Qo*Ξ2�R^K���C)G�N��O����pD.��+7��癯bz����V��e��W�H���υdդ���jE��8�@kM<$!�S02��M䐴����`��Q���c~ҵ}q0�^VN
�3y4
��n@���#�����=U![��#t�u�բ|.�o���>�kSd�����`�A3,�i�Ζ�V��c��%�6��K[��~<h�W@�#��T�iv+��;1�'DD82O����Ԓ�-`�r]��8l��U$�����ӱ2va'��]��Y��x�u��=K�k4����:�׭v�j��� �<�(h-P�.	�x*
.�42���;�\G�L���w��m취��\n���O��~�y��̞��<�����Z��������������g$=���Pط�#�	�ԗ&!g ��]�@x�6V��'(҃��+-�� ��V��� k@D�<p�DƁ  � ���U�!	/E��eD�ae2�E�6�H���7_Ÿ��;k©�4�����"z��xn3��B�V�,�ie��__��8���������wP�s��s���Q�c�'�aY���㤿Wخ��:�&�*,��]��U2\�V���~@b��Tu}L]�Th�F�w����B��W@��\�� ��T�1I������y=�ϰs��R\>B^^>F����I<�s�/�wȁ��Ŵ��[��*3B�BJ�0�C{$��/a�n�4��Ј����W����H�M축�z�h��,�l�9�1������i߱߼���%|{�
�ݥڭcֳ�q���B�;Zd�kE;���U�xN&����z�ݘ*vF�z��x(.=`l�\k��J���EK;[`��CG5&Q����G��>�]?VPR�^�-Ч��C�	Di�\f,���q�k[����i�͚�'�賈yCdne=�Y�(�apqU�Rt� /�F��v�e��"�qyC����K&E�l%�6?����0�wr�@�zg緁��|�Y�^D�i��X@�����P�E�M��u�~�֐]y�ez�b�4E����=.bX~aȡ!ZYix�N%�]���@���t
S�����G�Ɯ�n����4�Wu���~������ø�I�UM)s� 0z̐r�9�r
|H�[U$��b�N��*��L�!��v`0��.Tg�>m��chvq<3R�K����������=�F�F�D�[���ڣ<�?�R��U|7���K���o`�/���1��J�VY�k?�_GU-�h�Q	\����@:�r{>�]ݜ��og~�p%m	���5s�b9
�4� �ļb��&<vx��>�k��0��vMb<;P�l �5����$��y�P�3���9�j(�W�Re�q#q@�3s��8������{�:/��cyd�+xq`"��{��T�����O�$M�5�~�'��N��,��2��my�,�FMT'����5���o�3d�&��AOk�ߝ:|�F/����4� snQ�I$0Q4b�&,U�����c�*sͽ���X�1��e�Ë�J�%EӜ3@�&�
q�ղ�vc�q�۲������Ea��+#�e��u�A�{���[���P7 B�0������|s1!��s��
6���S�rz��Y��2�c��M2#N�z_�0��N;h/��F�>   � ��u�!U��v�i����R�'�0�S�Z����������2GN���o�5����A\w��#�