T:�sRX$�/�ύ��)�I9��ڈ�1v�W�����@(��d��3�O�Ax��/�8�gb`;)�a�bPs�5YUD��}��y(���ç���$��J�u[��7T> �u����S�4�~�E��"�a�m.�E3*R�ƉHLs�B��.�s66�Co0o�R�c|C  F�v��yc�½�pi{�_8�V4�D��OTT��@]����w��� ��OL=�W��]�R����ҳ�7S,y�qm#,b�� _kIy�+*�"�����:m��a�ǩq��<�A�c��j���T��IQJ�|]���es�74Y�	��~�X�Y]��B?���T를��D�Tɰ���s ��l�o��$��[��%��@���������(�+�����BG'[�xg��f{��0µ�dr��[4w��0�-�2|?��C�኱>m;C[��f�.}�;�߅˺�k�P,<`#��־�}%��"4:U����e��6+�;��،)��)��TZ9��QE�r1^���V���hN ! ��,��~{�pU�h�l��޷86p��P�J8��  
0��'R��c�Mm� �c`�=���U�ݖm̚ <��r�_8����ga�(��E��L��+��q��FB�� ��|�0����{ʾ!_�Z.��Jc�kz~(#w��I8���:_�?�G�!S V�l��{z�� -��<7N30O�,:,ⱁq���=2b�men�[��;Jқ�[z��Y�#6fxc7H��5�p����3��q/�D۫1�S*
4D캔�'�>B��1V�n���H��k�}FD
�tVo���'W����79}x�P$���ƆE$�L�����e�4&B��>*4�w�he�Hٳ���z4T&Mtۂh J��Y�r-��#BL���#�ThÑ���T
��}K�Vn�ۇp�w�Bx�3m �&f
���&��,�xw��a�#)�JL"Z�����Ȗ�_*v4�(��Zl�Ю�D
�ԧ
������*��������k�氏V�<;��0k�N��Na�7������W�i�ʸ�1�+�L)����Ԓ+!�ΡPB�ȽC�k�"�~G�2��>��v�e-�4�g�v}H���C(�C@l��
�|�=R*b��� o�Vbҁ��	��}�| �t�ZP������`{��k��XY~}�%��%������p�����3�$�jX�ō3s`p풓7����H��}�`A�v����﫰�Bsa�����.�.'��:���kQC�0����!Mø���1��|�F`��X h��#�`~��H�c�y洄�[��H� �62��$��u����!�'f(0��:��@%��&P�`�l����z$�����}B	y�u݁�i��տƞ�=�HF\w~�(�e0������U_�Bl~���k�<�B�Sy�!�a�<�Zw�y�m�u�����9.�P\����)wL�9�"N̷�����a��Ƕj��`��^-����7*­?B��+��z�Y��VϏ퍁���!굽_ʨ�Ǔ:��q�<�s�ST��R즩���2^q �������Y��vZ=����8Է�%�'T���͝��`���F��UX?d%�F�ڂ���k>����$V����s�q�CW�N����{A�[�(K_l�m���^ �@����Z�W���7RdX���L�O��k�N�<{�m�an��a����Ǜ���kKY� �rtY���oeg�oI�^���2*P˰0N��2 �u=��LK״u�d$aA��BJ�F%�!n��]��M�6���谗7<d3�D�3�=�yD��n&�ڈ������ ��w��s%�7�Y�D,*�4���g�e��g�2>
<5���4�Dy���=�v��D�-��!Î[�n�w�h|����F�B�2|��i��ASDy��HA�\Ө������wl�uh�!@�y���	���q����`���F0d-��t���uIr�b"q�p��þVml��V�˱Į&�7"�Ʃ��K0��|՟�eNY@=���d�(݆�>�X�<���b8p�X�m<:�S9Ɵ�7�O�cU\������iq{����ŷ
�{D:�/ݙ��Ku޼Ğ��}���|]��k»V `�aJ{3�<���R�4���*��8;�����$]dK����En!"�)S�5�����k�x�$��Cq�_��W5#�~�=I�-�no�vň9>�Q5.��gY��s��,�0��R��<�+3vA�g��`xŬE.�hC��W!q�W� �|$̗_���&gk݃�	 !~���S�9a=���O��_�6'��VL;:>��^GQ+����D\I���y�a/�<�I{Scr�%ɨ��|���ʖS�i0f%/@d���3�G�E�q�:σ�V����H�=��o7���������r%�|��qi�����Eܑ��a�I_����'��dZA�/RѻyXWJ��D��¼?��nO��o�;Tx�%�k(��;)(k�Зp�����KAm���q7��:�89:����;�&��͜W?�u7D��@��6qI3����Z4���Ź*!D�#�?5/�y��o}K%���₡��g\VIi	��F��6Q�+�m,�2�~�r.I�o�R(��º�P�6�{��#�O�=e�
Z��qg3��,7�f_��-�����G��F�	˪	�7}���-|$�|ޛQKZ��]a5�ѻ5�e�|��H_(~�-�KǏLz��^�"��\�E���L�ک�sB�	����4Lyx�0�gG���0�'�J���H��WN���a��nh7oe)A (�����Y��U��rqT>l�&si�)+�x