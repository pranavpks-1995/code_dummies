�K�BE�Z7�o���sm�+�SF��`�V�jN��9Хb�ʤ�FgT޺*[��4��E@	^�U�Ҽ��6���k竉r�(����IҦ��`�_�Z�R�Ƀc���&mVЪ&��1�4�]�H�Ob�.�+�b&���b�h���nh{,�8�Ԗ4��.���(�d�v�-��M4�����oqj�-ݫ�p�U��ϏlԬ/����o�hL}��UsP&W
�,�SN����bW , �¬[�����4_0-�ˮ���Jv�&��&j��i/��� ��۠T��S�nX.��>k��z���c>�!�R��������M�)D��Jd�D|�ً�5$�U��[����Μ�똔���4|�z������*>�]R�D�:��ߩj8�����y�qYN��{�M�3K��hN����q"�ib񒒙��W-�6q{nH�Y����s�e�%Tnn������ᇢq�(hD���=�����3��a���*D��r1�uD�N�c�pe�ٙ�5�׭w�5�cq��l�q2�<��P*��-c�q���-ǟrJ�YN9-�"����(w��]�6uY�/���Wwڞ���k���̅�m� ����F/�:��R#ۢ����_'�E���`ky.��4K=~��4l3/�v�e	�f��k����|%e�8; xU`�FV��S>�����ܕk�z�n'�\`�|5��ω�t8�ۢ��tC慍)���ͥ&�5� �������$K%���0e�J�𘜣:Zl ��_%dg)�Rg_L���
�� :z�&�5)z�ܥ�N�	�K����啎������$�+�B"݊��)HApw��L��o)���I���2)���9觡�+����^a��y��r�m,0˧��q�sߗ^����+���%����1g�-9ڰ����;~O�H�L�����C��]�w��[���h�ev�~	�Ƥ��'��Ԥ3�A���k���Z���`��\��[�a� 2%$D�
~����2�TxT�Xb[ޛ���p�`�7 �`Ut���V����Mh��m�h/�S��:
�_7���~V=%}2f��-���^ݩc����S[L���/ޕ�n�qޱ�5n���N-�aW0���2�>e���[O�d�����ʓ��3Ŕ�M>C�滀]�n1vU�0H}%�w�����{n�AUqYJ��ҟ�_�Yo*�����{O� Vq�$5; )�o��*&�n~�N_���Ř�G�3�K��\ih� �u|`Yu���E�H����� �ȸ�����E���㴮����	�J�vsLd$�G�!Ť��^�{@"��3��N�-�:%�R����o�"�e~ܣ�~��P\`3��EQA3���BLS��{�<hۍ��x�U������|KŀC�)���Q{ef�a�ٖ�C�[�jr���\�&�!73Z�cb��_b>N���ni\�����\�
���2_�a�j��7���kk�񩞓ߏ��mc�m�`�;v�2�B�e��R�����''�q�2%��+�?�w8k�"ŏQ�{�
w�,��T������*5/�y�Ifx��Ũl� )yq���e4�^���t��~2L7~��x���ڵN+��T�� 2��۞�Dgl[�\i�-?ܪ���V���
Nm'eXJiw�N�� ����#���GSP	.�M;g<�Z�a�)�~E/������9�eP)9��s=����Jn\���`F�X�A[:Y&4���*�CB�]Z���ujYFר_��SR��"��_���i���e���(���~��9s�>V�t���