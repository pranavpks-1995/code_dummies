�b0�b�jA���.��"��Yڦ�����Xt	8J�f��C=���Om{k;���[y��{(��W��;dD�@�]��J���iȔE���[׀8[�;�~	�P�I��ƕ?����'��>��x5ɼ�T������dR�y0�1�u3���t��T+�[j����g`��ߚ�-Z��cd�ä���_���(��?����	��}�!8V3��)CuG�:"�.�M;/G"F:MhXgZ:��� m�\�H�J�$  	��"'R��c�����M^S�������ĉ� �CFz�Q�B��d�nl �ݷ����y�/��Rzp�����UEp�̽6�M�ռ��q�����s���#����u���P Ѩn��-w���"M^~T*YD���%s$D�C�0���)�~7$���c���[B�x�v�G��v�Ђ�n�u�PEl���.��*\>��gg������-����A^��e)us�"kD��P�L�6"��m��Wm2����Ɏ�3��3�d�} ބš�K/�lY�Iw*5�����D�G0J�?����6=m.[�<��	iY���çK@�!z�O�:�j��5F8.M$(�ҝ�����$R#��s�c�L�
yiNvf�,yJ�0i��{��b}MZ���G�t��E�C2�����y��V���7+����Ҙ���2�˃��>�Թwe.4��:g�6
VU�b~= �'�Bs@J%/�;�JO����l>����f�������c��w[�9�=���@����BO���a��H�Oƙ��>��cX�I��J�Ą��X��+:I��]�x춱s9ł<�G"�f��@F\t���Kܚ�����e*��[��!1Y.䯶čOPL�"S\v���ai}���bR��}i6
��&]2C�[>AYsfS`n�h8���Z�}�9�c*�� ����������c�؜(*Q<R=_����tX�`�HS�X`�[�Ȝ����{�aP���cq��C6Hs�N
!��G6��e��A^��م�V���]�V8��>٢t`�4������W�-�;o�,��\&}`��C�rݍY�M�f�S�>�ë����E��JU�wh]�
�F�Hv��W���� ~��e;�<v��E��٤  W��3AbF�31����x\N�k5r���P����%�b�ʼb8wz���X��9Z�!��A� ��u�ƘV豌����*ĉ��U<C�حd_�Ӫ-���=��GBd�1DEC��v�ss�~�Ǧ���@�i��h.>)�.�J�.4���dŻ�^�f�d=����D�b�<���)����㴢�	���ے��~�M%�e]�e��{Ư'���r��u��:�(xV:n�����<���d����%��M^����t��e����q�l�Sw8v�x'��=���Z��ȶ�=jZf�m�7�-��ɕ�a��q©(�-9�z�,����7�!�h
�ؖJPD�"TVD�(U�Slv8*R.��!Z;{����!i3a�U�W/�2�H�������W��Vn��cM$��󄰊�.�k*JR��uI&2�4��Y��pwB��o�l7��:\rI��CO��tGj��KR���Wf�E����rD��� ���&�\�Q���c�d�:Z�F}�ӷ}97O��i�6���*��������(���9�B�Mݯ���d�^�-��+���a�mKJF��W_^�A�<�Ո�}�t�bV1"��gv��H68�펞h�ܟ���O���
q؏�PO���lã`�]ί��IJ2�3�M�AS�*6/�����J��zP%��d��/Z�w�*��%�%6�� l�5g���ki��������}�hz�^��%A��\�[�C(p�ί�����r?��:ȶ8z�cL�f��D���G�Xe�8��n4V_\E.�m^R��_W��+�  ���F�Cn �H������԰)�6�4��x+o>뻅#��w�Һ�@�R�_�c_'s�M�ǵ��T~6�I�>}�Bc�&jk�ձDn,�|���-|�$��uZ���S��VQW���Cl������W��U)���b�z����R@��f~��0B�i[�����n/Qղc[�x�[�k4��]�$9�2-�B��*G�Hg|0\��!�LMI���x��at�ܿ�2��
�`�+݂)5�?�
p���Mɋ���(����p�l�E��QA<�eT�
���)����>�1���C�7ЩD�Q���@�n|��ds\z����6s?=�EȜ��a����4�0�XaYѹKV��ע�K����+ezi��"(T���|>��.��3���?!��ʏ6��l��ů�|�7�k��|V>^o��A� ���
�>>MPY���.�Awe�x�l@�&r`�BL3u��6�<x>���5��$�0K����INW�fg�
c*��QX�&E*�m��<����6xpk�_�z�M	j�8~m$H�97RIC4.a�\�|/��v�e	�[H!��'a~�]+��_�ZX'g�'YK�l�kh��톘���Q����sER��j0�V�3�쐩TE��,��Ѓs�7s(���h��R	��vq�'����lJ[�P��wT�a���ϹlZ��Q�V�>��S���;ّ�
1�P�,	` 4�Ժښv,'��?���82��t���qm�H�z�����>� *�Q�yol���X@��Yc S[k�����Y�����
H�FX� �  P ���U�&
�]�e�Q��A@�)F�}��e=�7U0�C��o�j��\'z����R�e��%�JSm7%eN��J�>aC� ���C�X"̷�7k��e[#B	�."�P��'�X��I!��B��k[�I��AV���ɫ;��t�K��1���|L��!1#F���&���6pv�5G��{Cj�z7�M��*�T��u��å<��Թr����|@������������$B-��]gQ{�C�:��9�LΧ���k��l;c�?�%�z���8dg�0�JY�+�z�n�fn�C�EO���7��%�w�E]O����Ջ.�W��vZj%!��Uޞ�g�٫�9�܆����
*����f:0�Aq���2�;4JP��\�d1=� ��K 87m�k�f&J%l�y�$�)���4T�Ko�,Ck�c�1T(�\�:���
2%�B��rb�{=��ȍ�)�D.��?�ce�`8frw�ap
�]en޺��:j���ac�� Ww�g.%�-r��1
�p[�=�ޫ��XTXW�0s��ѱ�3���a��c*Cx��AH�n�L@��q�e��co�<��X灢A�5�G*�◜^-4>������N� WȋzǨқ5��lo�ˮ����&0��m�M~�H��|�(j-؅�=@r�����r���(�V,ȥ�3΀��G��W�Pr3��~H!0Z)5$=t�j�6_A>��`h�*�po�@E㍹Hx��<�%�Ӊߔ����ז�l���J��N'Z.4sڗ�Mv��'�u���9��|F���CQ�.'AD���6�A9�pކ7��L�F�CFL=�~m���;ק�A.�E�MnBd�ZO>�
낆f76��Jv�y�04�3�����D�3�#\<^�J[�d�F*z������b1�$晃\��$��9К33���ܧjy�"�rN�������GU������%�ݑ�;;���n�#���MT�����`M+����(�ؖ	��-���9����5G�.;|G����'�9Xþ�7(|Ϭ�3�[t0���ϥ�D�1��"7����Z��rDm�K�l2�a�m>�k�d��\��.���N��$�`&�|�"��L������4�dXmYU�xQp��s��tV؉M>�>����C(:�� <��|Ȧπ��r_TH�����M����t;B|�N��}$�'���)d,w0}X��� v`E�-�O8�hA�ď�2�G�H��'�!�Mt���j<�}u��?=*|�j�'�	hS��d@݈��q�
 �g�kw��|��%�~�W�)ϧ�����4�S��δ���4 +�f^�l���އ��B�:��W�s�\4�:��MDSy�T���];�U#�}�U%�?U]1t�EY+  |xY>��Ҕ6>QW�x���/���b=<��9��o��#(�'�7d|���f+��f`���mL� ����N������R�lmܧ�a��>�kq����)0�,d�~�4ʒb��b�i����@� �g�d�hXYB��Ɋx���opG��.g��2G�^͜g�y3�	\@[-,�1��ٺ2�:0��O	��u�O���w�k\S��F�� �   � ��u�&)a�dba}&C@�BHw���Z��9�
�G=�cf�N#�	�@�@�e���ZA�c\�r�
���W���|�� �s%f�/<h�=Z�!�e3��Zh�Z�4�h���3��q��F*��p��4Iн8Γ ��#Mi�P6�C�E\��Aܣ�u�K@�q��@<�@�RD����l�s-s��l W��|@�{	��%Fl��	�i�/��5Q V㭗����F6[�a�� ��Χ��	�����!��Ұ��Nt�t�2moi�-k�����E�aJ�kt5� e��2�jK�*��"W�����Y�尘k₸�BDpث�_�#T�������kK��Ƭ&zpvX])_������bN>\���K���##��W?�|�ݕ`�d+���3�;�A*�r[:�4�s"�鎨c:*������:�ݠ��{��*�tV�N�W�TT����f���/�I��QI�E�~Z7�~���C��(�۶�⾲��1�+:2�4y�R��9M�J��5EJ�y>"Fuǲ^�*z��:o�	%�T��[}���LR@���;�a��Հ���@����"���P�=y8	̡��Q��r�����{���{�J��,'W�G�B��SѾی�Y�� �7b>D�� I׃*d:O���w���g��&RN����c�`��Α���)��i�E���يT��gj����^j��O�Xԫ$��)w�t��{C�[4�~���CY@��Y��"����N��xHm��DhQi�F[���
�D�MP[�7����5�y.Ӯ��ӂ[ݕ��K[�g"�&,�"�7$Bu��=�t��s{�ܐ.<�P#�S�R�*�'0����hLG�S2w����`iePmv1�P��	a��`ta9#�o,b4: �^������-�qh�ԑ��{f%��"oB/;͛�+ͰzQȇ7P����͊�>hsy���$DMĸ�v�F�)�qu��<�aV�`ܨp�VRP���%�Ҙ�Q�DgB��XQ *�=В2W���P�"2��Pxъ�e�����ZG�?%�0ߨy)N�8�q�ӷ��b����yF���z�"g��!�nf�b+��N6!fY���T��ηy�	3*��D NN(���7�v��	ƉC(�����<���P�@�p0��2̟�T��TA�x���j��E�rA���X��B�=N�P�0]�C[l�ܦ�(�s�@`��0�(h&�e[��'��T�y%�Qkp��N��Ų��Z;V~!Z��4C	h�R/�2����|7�='�2�g�����W������V�dz���F0����rK�qq戠�/(���'�5��^{�ǥ����r�X�e;;q�X8�#�]s*��U�P�� ����ٟb�p�6M���y��ہ��V�7��FS��F�ũ�x���@x*���魱����_?;=n������u�������z��,8�S��w�"g.[Ť�[�TѢ��U�0'8���&9=�/.�����!�v ,u������[���Y�\�ȷ0$�۸ _�c4Q��
�Gg\#\u�,H5K�u9)��Kl����q�1ҭ����p�b��Y$��5�t�"w%vp�s�U�����L�i~6�%�#��q�>Y6�gm��;�]���uv9�p?W8�D��N   � �B-����9S]	����c���`��Ri�J��c�xh�2�NR�託�%��RCgAz�p��i�D�����G+�1����0ǣ�w}�|X�u8y�dPY����m���xȞ����r�tzVH��ԃ	�~�: