��\.�Jc?~���މ7����U����C!���I�5ĩ�������$�� �N6c������L�|���8�U��#9�@�˗��>	��p������̕k"p)���E�����K��jL��Iz���_����z��A�?P�y �6��!+�M_v<d��ɃzI� w��0���҇6���Y��"�d��9(����1�$9���H���m��_�F%u�B.���vI��`��cV8��e��DP��8E�h�:�ϔ��?G.�u��Oo#ۘ�A��+�/�m�c~����<F9G�Z�``P����O�w�̜�#��q;�b(.����� ���UG�5�{ ��{�2�Qeg>έz
��զ�7�p� B��v���g�P�%�Yf<����&�ힵD���m:��[�����lVA��%W�1)x~���z����W8H"�=9�+�C��>�;Azs�~,�!�sDZE�8]�>�˿������X���(����X�PI5�,{�6>кr��@�Yj� ��,�_ĸ��9v�Qy:IG�a\��R\����E=n�5��	-^$�a�WZ].�̺�����y`eS�>��je	����n�'uF?�]'w8�'LY:�?A7��Y��\4AnC���l�Y�.�w��D��M
B|g��:�U��x)��&^������x��)�#��5/Ζ���i�茂+o�r��