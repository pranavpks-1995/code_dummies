�6��iQd_	j��ff�����Lp�QhfI�/2�u�k�gf�W�o=e�w����
�yq��ą��)U�3>'���a����<�ԟ�S�c
(ZV���]u�;ڣ�ɳ�2�)\��zw��_�=�䰴�l;=Vx\�w�U��9�lX���/Xj{_��ߪ�ɹf��F���
�ƤZڣ���Fɍ����k��@(>��[jѺC���GZ`N� m����� @e��%�Ó����~�~���fB�)};�#�-pp�P共��x� ]q~��[��rAx�`�r�B�g	�2nT՛���_$�[Y�������̦t]���\��r�ӯܡ:u�s��4��F�J�5��� /#cD�	����F��53%
�N��l��ƀn[Ƒ�Ɲ<~�Kb�@h`����#�Sյˑ�T(��u1���QЃ��&5�����S��7�=���i;P� -��C�pJ{h�dxx�ӷ(�wy�m�H����T {1z�O3VU�?�˝h���qr�h3W<�<��LJ��)8ϤdѺOT�R�Q��x������>A���g�K߸�n��Ʌ��m�C���~ubA����ρ��[��x*0E��h�FhL�Az�� �I���i������S4T���K�E��#irǍ�h�1X�wV�e�Z_l����T@JU�8I�焤�>�0JT�ۡ�����M[��M�l��_]�����0����U��C#����=&�򲷔WC<tJ@`��+�y�N�6��f�X�D�]�`�h/ۋx=�d_!�7�~�Q��<*>�F�-s��m��O���&�Ѵ��-���6����{^��1����k[��D�OP�h J?�p[Zo�\d�Ȗ�t��mk���^�s����BL�x����'6X�Y�d�n&�7LaƑȰ
�U\v7�/�l��j���Lȯh�_��w� �����|ầ�#+ʕ���]��x�t�Ce$@k>3��f�Ddv,�����9�ɥi�j(����ô�.�t��� #gx���ܺF!�r��5���yC��@�6_��ՋƠ�%ʗ�ӡ�n0���=^����ؚ�4!�/�v�'>�u�Й���o���kv�Z0glV�a�x*�DY�H�"|�6N��;ɬ��F������\h%��!�"y`��ץ�J87J��$<Σ�}��i���j����>�]Ё�z�~X�M˚�Ŀ4�XV_�l�����]�$=|uţɧ��˶���[ܴ~xm F޶n:���ŋ���̿s���B����Q��a�������X���l�PU�Hh�y�Ó���K]���
�PB`��e�����g7�D�7bmK2�WE�^�mcⱓ��K�:|��
�w�;\�0vg"16
 ��h �a� 2�nsr�Kg��H43220�1u�@��RD!��rU��v�7$Δ�z�x�-F+�W
]|�ESlr��6�Z�xҽ����F&�8����F��G"�T   �F�U�$!.���R�]��<C�\H��̃�����h�I���@<����,J��Y���C�����?_)�Y����Bb��X5R[\��Z�4�Y�/~Q�I���U���-�G;`���Xi���EԿ5�K�o��fI]x��zx��O���k"�N >��4[x�t�88]����l�_��KA#5����v}�d�!@�v�4����N�<*���y�R���t���v�gr��<��[UHa5�rhE@������J��X��S[�c��rħ�����h~���Xt̕zz�Ox�ȯ��;�|J\�=��0�Jދ�-?�4Ī��QZ�P�]\Q%
���_l��w"ey����(��G㐨mE�{f�	���`��	rΔ�Ք��1�I8�R�Ļ��cG"*F��;U�%�[��9����#�N(�6�����扫6���f�c3�a�b�3\�s��5}tAz5���y_6�vvlQ��b}�q�X�x�:����tvJ���[�w����4~0�A�i�2l���+���/I�*4 UC�S��f�����%اAp�4h�zF�&�렟^K�'p��¾mhLU�dK. �%��/:lD���?A��*�F����z*y{2c1Sз���>3@�b,ԓ��Ud��/7u�dz8�g\�X�&��y}�i�?P��cg$s(\��gj�*?.X@q��5���n�H�I��4ı�%����ϙ�w��z�����y�j�}�-�,�V@�&#S�!�� ���tM6����_' ���	~1�]c��c�s6|��~���O�$Ì (DM��?ά�l&`�DP��	J��xN��!�&9v��z����lu��?�L��x��h�O�b�7�J��K�w}!��i��7��S0����?�q��D�%�χ�--hI1-���U|� ���0B���D��C�fҦ���y<F�@�,��:a�]a�a��që����(��9�LS�!����"���Т�J¯��r���Ď*;7��ҳ/�T�W����5�ˏ��'f%�%zwXғ�������>9m�L�,%�yE����84��qX4��� ,�^���!���G�x������8�u}��`�2Ud���7׬[�9��_�����:��_c�T�f8�[�p���1���|����������]ĄPz����bo&��@�A�����v��˂�>������oY\���V�Ǡ��/������&Ǥj�*��lp�<d"dU;�f=�tNʻJi�.��.�VI  S��vd������ŭԯ<�<� �F#h��PB��̘|1�	{c ��!-�Y>F���*��U�N(�nϿ��,�|p$����p9��%mD�����ҥ�ғ�ԏ�-��	Z�o�ĮH2!��lZ'��l�4VU��ZZ�����T���;|�Z��dR(��.�2�ٮ�F}�cruV���o�ZS�����S���w�5ݗMV]W�.W��Pk�;�b�CǱ$.[�&�u�ɵ#�gI��XJ�s�K�Ao$�a���j��^��S�{Z�%���)!]��u@"�*�K+����0��+U2�7@�V�&={����K�Ҷ!�)U䡙;�OXpu�L�-9s`����R�rk���%�ej��N�B{�7�rZo�s����<�N/� �p	i�p��� H:r�1D�W��>�z��2�'gM�Y�q�R����Mm ���O���}��`m�������!��W�*�.�o,M�;��ّ+��p��0�GN�~   F �f�u�$2)-K)�����@r�J�����	�	V����� ��ñ����3�9��Uh����{۶�l:P	�!�D�=�S~����f��,2	����t[�	��O���B���&���� ���`�_�v�\�:�Up\
]m��0��~L՚F��n��_�Y�?z���Q���<ѧ7�[}�%�r=�|�����n�4���������t0�	*��a�����q�uF�Dm�(_w"�h�s `n��B��N�`l��8 �wD`��ՈXcR1�3�D�PW+gɝ�1JJ�#cgu���SN�w:څ<j��7B��v��8,jKcQ�V}:KP�n�Xx��1s�p���X�If�[=ۼa�z�9 iP|
G8���h��|(���aX+���?�03��`�
�|��W+ NL�,���IR�e�٦EE�h�2�[��N�p}ͧz2S���\�9��+$̬�,�*����u�8u*�	c�����`/�`����P����Ty{S�6�A�uk9�8�/[}���
v��d�����M�Q�R��(DQ�7��l�m֞�R&�_�EQ�\���y�_�B�����6�0�� V�QA$�!�y�M�S�:o��C��Y������Ѝ�JK4;�3���v%��2Mo^1=�BI��y�M5c�/X����}uI�ս���/������lUf#���M���z���+^�߂b������v9��hQ�"��� 5�o��15,5D�.A�G*�UvI����H:]���G�M�l�{i6�4oA�[�g3ڊBhX�o#�fT�68p��k�c��THXʇ�I0��	f,H[�i�D��g�q�6��q?!Pq��cEx�vH�F����VYZ�|n��c����Ц�])��E� ����T�����}������V�HE�n����js�O
��2뮸�B|H�C�,<xa�+�T�5��q��X�*Qɍ��g�*��	�wM6m��j��~�h��My$�k.H���LV"��{��hvw�1˄12ؕ�=��L����U��I�µ!�P�)�5ɀ�6��P�M,��.��2���p�b���0�|e������M��6V/��v��J�C�����ip"Sڞ���j�)�P��D�f8T��lzoE�Gi\�\y��?Js�C�Ê��?�hkȣ��M�Սc8�3�k��5M���+��s���jXVOP�a^�3ۭ6��oS9�z���m���enė��!p���m$_w�� ���9���)�"���q�Zcl%w�0u,���y�Q�3%�@dw!m��
�cG���=�ÔQ�/gBK ���:�g#}��+� v/��~8A�h��?��@j8��b�Cx��Ō*o���1UX�������G��iz,����@F5�]����+����Ê�_;}=V�E�c.3M�l2�?�И@��H1��������4��i5�We��I�@)�%�̇b��O��@���U�m�C߳�>_�aF8+v�b�o�o��;�z")�j�5�d�p��p47�)ì�N��{�J�ja�4b1����pKFaG^'VǷ~&	���g4]Y�����=�kʣ�:%�q/�G�N}q{,+"p���
%�?�i���sS����?���CIfi�L��a4�=������f[�^�H`Bk8����(�Z�K���Ŏ,��9��ި7L
��MNr�i�� _���3��:����^��WT	4�,�+~�z��e�|�s+�ԉ�ɽ!,��pSB�x�V@e�n��ьo� �v�7ƭ\�:k^����5��q�(�[�J�y�r�