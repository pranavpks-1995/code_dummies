.H�D����P����ʁ��$2� {fW��H�d�B�Fr4�����������
��>Z��e�3ם;3\�:Y��筿%�e�Q'���
�H�Z��Fj�_år��`��ׯ�c��B�Z��mp�� �����_銫��TA���-����
��v.r� �`�� �2���p^JV?�#���� ���5uט2�H��!CI��ɓ��_��zP͇��J#��c��y��F���6)G�))fV�J�ނ�矸e���H4w�ExA!��p���*YBk�Y]���j0���srZu[5�i�q��>� ����t���[8��#��ϙ �/��5`�b�y$lF2��"(���Y�,n��磙���.����|�d�ᰟ�m�M��5bb�5��+6���|��|����9f�?5��]S���&6���T��Y��q|��=u��Z���OS��	��G�F޾��I����"߭Ӛ)QrY��*��km����WO�E��_���}SҎ���*�fz���J�!$���}zC"a�K�/
�I
��h?flm�����F�]���C�yQ[�t���&�؋h-@K�E�/��v�a2Ro������5*��L<2P�~)��~�A��W	F5��6�}�^[sc�c�;o$S���%��YӔ�LW�d'L�bu, F�H�[�e�B\l?\��i	��6L�{Y�)o� �.�.}��9����/qW�yU<[Џ��ԨB����5�.�5���̋.Dv�B�Υ��.�C�Tvq1c�Yr{sm|�P�O̾�,���͹�:o�a�,%��8�����W�f��|PC���_F�;n�r�e6�r	.r�{����(eC���l� 0��I}��K���� WG9�i�G��l��ڌ:ƫ�V�X��A����@��O��w�J���B���)�wܴ$���6B�[q)D��O��k���8����V~P��x��+:E�rZTb�xɊb�=������ݒ�=W�":|x�n�j�r\�^U�z�sb���9�l�Z��}��yG�5��RU\�0��c����F���p{�Y�h>� G/���o�>���ȹ^_w�+�|�_���]�B���)��(�9?�Ze���a#)�ʴ�o�v�y
h^����T	@G�,5��V���hY���8�&hK^� }%2ϟ�,�ri����b�\ �W-����.�Z�r<�����"Sk��5�W���0�oシ�=�0kO/S�+�TT[��̗��3��g��\ę�D��7κH�c3U�iB���{%(!������` �EG&"�s���N<���=A�e��8Ip�IG�KJEVu�P��%8_hq�C�fo�K܂�8	�d�eVX����՜dg0���"� U�#G���"rC+ �|���
���_ޒSRǂ�[L6	��6ņ�t�a�����b�4�V~P'�=��,�"E?���Ώ�¨&:���ģ�WQ�2ySԊ���Z9[k�A���lxs@Ӝʎ>)6̇�	-�,��jIW��u�	*���� %���b#D����a�IWˋ���$�ޔ�J�]'��QF�NV���$pJ�-zĞȜ��f"���02���<5�P�mq��7ҳ��%�������Z�Xƍ�lޜ4��y�Y�.���uj�dM�:��|�'4�-�|��$��p��m���?=I�ǿ�/E��C�8r��z�J@��W!��e@�F:}h��0�jt@�.EtW9M݈P�-��R�k�Xä���l� ۑׂ�՚��0� 'z��y����Ԅ�Ъ��f���_J:���S��՟��Ȅ+��Zf!¬0��bT�f���.�o>���%58��U�� q��8p�Q�޾ƣ���ȼ�\�H�9�0����ޏIGҶ��8*`�j��Y����(r&��k�\�����z;<Q�wiB*Ȼ&���~������۠d��W�=2��^����y�E�.�@�\�)���Cc���y�f��9��p��Auɾ~m�����!M�m߆��=Ҷ�@��p�ڌ�ci�>�����4VЇ��7��s8w>sp���{��$m"�|{�-g/WU (~�J�xy�2����vz�>���5t0ξ��B� �Pin��!J��h��(���㥲X)8��{]ξ�l<�n�h�̰Y�=�(�m���W�.A�D}�E'�k����Z{�_�]Q����|d+�g+��~h�i�A)��B^}�m�!�rk�	��>���������}	%Bf#�J���%O,QR[�e<Tnҭa%�c�};O5ĺW���o�h���������3�og���q,[{fwN�EK&O5�����A�A�� ��Ǫ�Cf�֘X}�f��� ��w��F�G%��D���n��i�}9�C�H�x��!4����}�nC�t���%zV8\���nx�fi��.�3�����6�Қ��Y
��6;
��6�(�w�^�>��GewB�c�����t{=N�$I���T���,q~̗U���=�g��e��&��S8Y2��4�h�v�0������%����?��]�M����D+B�4�~��h.s-X��~��%��j7�������o�!��C2�X׶��k���|���a��}z��.�"�_�!��5L@d[.�.�N-xS�1d��u��	g3ښ/'�{ϒ�f*I�j�I}귚ƒ�m��HzY�y���M}1ޢ(AL#�`�+��?�J����	<�{F�d��#��m�W)H)��f��f2����&�D�;�1R*��$/�67�e������d3Z�M�Y�/��0�^;�n�^�T�����'��_dΔ�{�l�j�Đ������F}*2��*�� 9V�O��PH�8b�0\�2�Eku�?�	���N�x�>�T���rz?�Zl&;@���0C;���I]�[`�/�H���� u�3�t"|�}q]ޕ2em�yIq�L): �l4�%���2������й2c���t'H>hB�FbH2��Gʤ�T���L���r���W��?�Q�ȇM��'����8_j�Ű�HSI �i����M)*�-����,��^z	��|ą}���1S�%/�4���2!����0Q9�1Vyb j�tz�F��;ԑ*��T�T����h��l�35ym*���Q�C���S�[� ����<�s��e�/c�1f��E��
�\ߞ��eL���/9�lH�@�mxE��ezݢx���0G}��u�ڕ���U]b�3��5Z����!V+}��R�'��Pt��jW�u&��OlL��ٔ�21�c7�vC���g;�����8�1uUz�6��P��i���c9ш0|�*�	����-���x����5��%��C ,��t �{l����.uz��t�3A��%%u�n_&��5 ����1T��W������h_���nH�u�#�#�ei��[8ֿqı:�.�����ך3|����x���NL�/��X���vS��~!�m����-_M��oLT2�|R+el[���i���C/�S�߈��JYiu�(z,�7���"������[� AC�,x��]	�6F��Tq����j�Yci�Yt0�ZͶj
-��f��Io�ѓK�C<#������6���?���i�B���}0����Yb�����$ѩ�*�wn�^�&�e�y/�eh�*�6���oJ��(>lW������h�W{�n�G���L���MG�N�4Z�����)�f_�N�v����hw�0�4}F ���NȺ�rx��|ʍ/\���?%�J��Q�J�0$G��i9J��B2�>2,4 T����g�x�L�-�(5*���흞Z1PŸ���g�������e�U����%�- �s6JXf�\��5�/o؜ͱ���g�/�mM����o���xQ8v�.�c�6�|Qvb����B�`z�O~܋䩞"�$G!��|��g����C�h��j �?	i�J��q����Z,� ��b�~����^�=blV�@��ӎ�~��r:���"�4�.5�W#x`h}D_W60텸`�]�nx�!1��3*����l���;��4�zbĭ@gbt�-�;pՂF��Ŏ��$�{�����U�:��L�wL+�T��E�΍.�0	d��;)�E��xk%����ԑ�u�t�x)mj�)ZI�9��Ƈ��~ıw"N��j3ԭ�ROr1a���яy��z���t�5ս�S�t� ������>�Tk�]�6��}���$W�E�5�SJ&��ο��(���^r
�=�����f��0�(��.��X���H�YW�(r�E���Y[K���/f�2.��[���Q�S]��#��"�a�3��ȶ�y�:�����7�vbՐ���W)������ �*�h� $C��a�l#B<d����
�S�X������V��J�/���y� ���>3e�Z�`���!��T�X����la�D; 2��f�XI���w̑>O>Ӎa�r�%XIc�moښ4�L/!���e\�9��B3�Q�f�;���	��б2�@���^�k�'�nK�G�Ґ"�m̹Aô��T���np�H�H�z��A�%F��6� ~�$�� �����"R�S��[av���l���ݧK۵�'�1f����2�'П�=D����>F�Y��f���
ؙd��������M�J�]^���!��3�ʅ��At�hKN �	Ќ]��Y4�вT�/�.w�!1YBR<dIU��^���
�����R6yN�Ŀ۱�\�0�(e��k#!�uJJ�D��C���w���(��B���`C(�9�@�����'����e���J�u9(�!u�灪z$w�T��Ch�)�Y����k���$��ތU����0��U��c;	�T&K����ȻI>e�~".Ά��h�Җ�v$�����lD�����*��|9Un�ƽ�"� r�8�s��D��������ǃ��4� Ex_pf�R�s1�7
�޺~�}��X���HQ�34L\�=.k�yw
��� *��ti�yg�H��I�T��Su�1�;�ӳ��"7�(ʀ�0*]x�|I!�Ԕ�5 ;&oK-���2�++��^5� ��1��<�4�	>>5&���� u���&�Y�0G�o�s��N齿A6޶[�9~/�ȇG.w�,��oԛ[e#�I�t�OT:���k���+d'�U�s:Q|�[��W�=
��}�����
]m����fݧzM�>����fC�"7�.|w��p����k��4br�jPB��=�q?|b<",��H'yk�����@5�9�do�O���՚��h���t�(؟�r��|<��3�m{�1&�u)���d��0p����Q�"ڵ>���8�y&�N��
3|���h�C\��ǚZ.o�R1��r��9~�@���Otm�ZG��G^�9��G?���0��D��.�dܷl�,(��U[Ǵp�Љ��^�:\!d���7i�y>͂Vw,�%��b0;�G����0�n'�AeДkh��p���T)������%d��s#;�`��2]*�c�
6?2��[�� ^!ޑ�a�wx�s�$��'a��J~�?��E�#�=�H����W𭌦W;qG��uį�]d�d�%�/�Y7�6�)E�V �Lժ'ϕ`/~D�a8���0��Mm�\����A�Uڽ\��!4�qor��dRS�K�t��zh���񜇘����G�5��1ec��X���}�[������Ϲ܊�S.5�T*���h)k`#�^P	�ϝs�ZcN�;�;��l��#QmJ��>=�Z�o-U4�odz��iI%~�ƒ�|����#,����ln&+�ǳό�K�Z��]��L�y ��rҕ�"����!~��i�M��>�>Φ6�~��oNx
���@�(�1w�'�Kw���>���m��6���V�Cqf-`&/�h2���z�+�;���Ჴ邮�$٣Uʩg��T��rƒ~�~�T��R 9��I=�*!���k ��a�M���y?Ӎ�Σ�Z�:���XQ�NBS�����8���n��+�� ^�)�ZDB����"Z�~�����׌�������s���&�^U��Đ]���qR���ٵ��P���Z�߀b�}9��*�	"
���DlO���|������RtS��{�G"J��r����S�+��L�A^-�����ϾU�I�ĒA7�n�%�/V��a����@A��?��~��