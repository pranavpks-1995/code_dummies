��Pt�����`��3�!�1-�&8���(�9#� �Β�"��w�w3
���ę�	�Bd,,��nJ�\k-m=��B��ZM;�m���n�ɯ����]�z��CʽH�h�ֱ(�#�_OY27���É(�������IM�V����n��[��j	�q�
1�ko�`K@�b��${a��?"(:��W��S�X|�l�[f�3 ���E*��d��X�,~���-����ၐō�g������}O���0e3��v�.���V@�^�8<r�	R�p����A�����Z��BO٣XС���UpU%� �_����fu��9F���-���$���G�s���It��U�A�
ϭ��}�Xe4�?fX���c����hT��q�zS��I�.�9�}{�� ��S�C�����$A}�q�����3������^^ �8n�5�^u#:�hei�dL���YU{������7�g"}�Vp2��)�V�+�ﻯ�	����;��A��RFh����~(g,j�Z1��C���v���3�,���H��TQ�p~���Fx"�ܝ�A����0�5��L#�N�� �ˊ%q���6��o�4[][�4=��`Q�J����G	�=��P��~��I&xI����hd��%�3nh?�wӨ���-�:z�\d	s��y��iŐ�X���Hs�i�^�g��vo�8PN����K�LA�+%�pX%��"�7��e䀀�P&�wY���!P&���&�l�B�Loi{\A�щߩĕ��<��m�l��Ͷ`Q�INN0���O9�^V�b'y2����emOh�(�7���Rש{N�\���x��%�}���W|�![ǃ�.�kEJO�+�j�G�QB��4:G1�x�+��|ȹ�ƩJ�����|����6������y|��\f/@s��b7���'�V�zw��h[�u�X��"��Ay��	�N���:\?7���Yb�o��ТzU�Qq�#$~��p6���\�*�n�`�B�v}��߲�d�eg�A��o��-jFb���d�>�Ѭ�E[�-e��M�-�8Ց��s�-kc�˲��,�I�]T�P@�4Vi��� >���D/b �����&��?y�g�q(%#�ϒg��������