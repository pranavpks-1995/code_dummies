��`4[e�%�S�w�j�ۈwirY�u&m�����}��JƳ�,4|�{�����,:-\,��1�z�@���pUwP^%$����K���Ȧ��i>�vg��� ���HA@���U�xM��m1ᛘ�`}�D8�F���eG�H ���~}n%Xi[v7�AV�X@��G2������w.	5�ג	�-n��e�����z���[�Ѣ��Ip�X`x�|���i	���$�6����Nl:�Hm�`}�)e�w�����S�E�,�	����	1�e�Z�j[��%+~���M��z!�V �
���q�>�6ϡ^,[l�1��Iz�oD8Z�rx{{R�݄<<0j�\� �����������~�Um_��ڤf�Vڐ����O���X�b�-�.����
&�,�mY�����.����j�W��C���
����L������k�q�.��Jn��X@�Y�x�I�9�,��1(_�j~Ӎ-H��F�����%�m@�|��RG|�2���h��	����?d�u���h�Bs
7�XU��D5J�ż ,q����gv��@��P��4w�UyR�"�/�_�;�]6�8�3���,���b~����o+Ue����1n�Z���Qf�Z���T�=�M�bU����{q�\�?"	r�h9#4�p���Z�ټ�/@q�p1p�o
��F����������t�_;�%]Ț��M������rؙ�IىN���<I�_������n��q�W�^�"�V�+PA�ꯤ��g���ٮ��2��^�Y�%���!�`LjEإh��xt�?TE�%�Z��mS��fgлX���l�́}�Y�`�$�L�-Ɯ%��9��H��j�=���=��Ca�-�E5߲�د9
=w����+��J0�Z���g
��bTG/,� ��	�;:\~?^�	��S;g��B�����Ɂ�N�m�R��'֙eut�z�����88��پד���~���=#C�A�8�U��%��� ��ʛ�iu��m��z�0T]�P��m��F.�/*M���hFs�·Ut��^����z-*���V�G�T �Dԗ�����3��^�j)K�7�M�5���}f��w�k6��􄷋�3;�J��멝̂��˫�4Y>�X�َ��SGX8���[/R(ٜ�\]��mz��0�R��c�P����u��(�5�
�͢8��YB
��hV�-�:�A�����$��Q��\.�Noy[u=sQ��U��}F^���|�@;'��[6����L"b��g�#_�-�4RX�y���`���UQ�����zy#W��=ฉ*9%h^m�D^��   V ��-����a���l�}DR��>��$.�R��|e�b0�)3�[|��t��;P@kC�����
M�^��m >F2��m���Kxxv��J��>�Ho�ځo��@3C���Pj��=���]�%��o��ݣ%���-U��[*Z0w��-s~����cm�Q�Z0m��L��7x�'s�c!�,$�>��h�c`@oy�����u~�d���Ô�� ��WC�;tV3JXk���7�l��l�?�s�(d~����&�����{�i�� GbL�z�Ļ�r��y���IL��>S)�ڑ/��Z�M�k����V_��(�*]iSS4D�
-��D�����a���_�;U񈍱�|Q������؀wg��f����g����U�Խ�^�{�?@���$$�t+�D��M|:������WvQ�@�G\4W���s�8;���B-w������Z�	��U{Ӣ�Sm�fh����2��A�C��[�ߛn6[�׷��y��;:�[��4�j�Кu����ל�P�)�׻�*o�f��C+�pC�̋�Z�̥Q�G�ڂn����}U�!���Ё�4������+F�&�M�����@r �?���[�	�0۰C�4?�5	Z"����3蜒a�Et3��r\�@����[���I'��.����ܔ�c��&2�t�W��-s.�*B t1?z�
����� ��!�]�P�g��GGu�q��S�-�W�u1� P���F�1�P�A�@�����}�����:Z����"��U������ ��k}=&��5�1Ǒ��5t0�=�b��UoG�`�Y����	P*��E�� �l�Q�ھ�b��o!���ک$�W�>� 8Ӂ���p ��~���i�����Ku�[˜,�o��j�>Y�:\��!c91kR�o��f%��!f 
��rj���x)՟L\�~����SwP/�(�� ���'�ȑt��';+���v۲Ǖf�ڙ�W{O�*�}8�/G�' m;��9����g�ry�� �`�ٿ�&�@7H�yV|Yg�´��c�,�;���ŏ��̱Q�R��K�q]~��,>��b�)
$�msԃB{�E(�f��������!��*Kb���B�  A6L�b���&��~�/"���-'3FJ|&��Db� �Ji?�����և͑/-�?�tXRкFe^yϞ|g`�$��1�-��L�,+4'+�����a`XF��X '_�" Y���2 ���!� �o�7p��\���۾��X�`    �!��%�b0DT��h#�
��`��Bo��H�\���{b�U����s��<�,�;<m�D�?��z	�]��1��
��]>����\�c� ��՟��Q'�g�_��>��o�?�X