���H�4/̕��l�%ѻ[��|�'�#D! 5|�N�;�AY���.���)��zs��e���T��=��R�`*h�c��-�o��m�r/U��������~c���� 5�]�u�3�kO��y���Q���ҳu7/�\��h�������r$)��hﲛ�x��7Z�&},%�P#����hP��I���R&�}��Z����J�ѣ+�*m� �׫����s
u7���;W`Ѹ�d���3~��b>�Hp���X���`ey~R�`��g�ZhKǺ�-�5�Au�)��rEUc�?O�I��V�l�F�����c�����5S�-ta�0^O�3o��0�������k�����%���#�Y� ��y-�PD+��V��oOW���i��dovb^���P�pyw�a[S�G�޺�Ԡ.ٵ���}����X=����-��|�� c�rv|?�X�/!���{���K�s�ƙ��72��9�*vq�<|C�+9���]��K�+�V�׌���WX̊�&�u�����u�:4��dr�sڀa�V�zS������ǿl���[�!���rm4��}$#^V���:Q���}�/�'3�?���������i� ��4���
������B��)>�� E�U����D2#��w)�ڀ8SM t7�yW׿y���5��&Xc9d߻'��~*�E�Սa/�<��5rf�C)�85TS�3yO~2�@���C� �g%��f��Sm�'
�{w|3���U�؁r�YY0�v|	�휍��|�������[� ������w��7�&u���֩��ZX8F(9l�0��H�nPq8c6�0�uԥB#��ΐC9kh�zj>�Q��7=���z!?��Z�Q,|�+	$��~�;��4��<�o��U���9��p'��=F���gc��	�/���V��)��s6+*J�sU���W!1�$qF2͓�y�׷�ؿ���[�p�F)M��lT�`=����nD��`���!+
p��JQ�^{m�p� u�3�E�O���q�y���'�w�`[�};�,.#���b$�C�6�͆H�m�2�}8B\FL��c�%tU�5���׶�sV����$���D� ���7oa*"�|�������Vi(�&�������ӓ䎠˥�|���9�AJqf&�#��}�o �Ȩ����D�{��6�ri�MR��P�H����2t�,�"s�~��̲zi��eW�Σ�BO  q�Hj+`h�gg�s���M+��6�e��~�s�%70z^�@&�3g{uڵ�|��`�Y�T�܉��/��pij� �'���!V�Z �7��Ê'.}c�-��T�+�� J(�wP��%G\O���"ED�b�W��w0�k��B7�W��.w2KՇ