�]Hik�b\Z��%@���f ��������k2�1*"/�a?+Ңo�)����aOU�u�g�� ���ӱ�CB�� �Q⤫�����;v{,e`�,�Z���l-2�48삵D�	�-��!m�0z��'�Pq�d�$�٥AY���	�׍��Z�PO]�6@�Y���By�x^ՔJ��|���I
��6��j��`��%�!�-?�ԍ�a2ċ/u�Nm>x.�'>଒lCCS�=���ӿ�����}f�'�$�����8躪�웶�f��w���&<C�m�0)�f��C�\v��dV�J'i?Li2�B�L4o���1@ܫP�_�ֲ,)��p���o.��&�����6����~u�&�V��U6��}�:�����a�4�P2?��(�s�AP�~2��Sa�Wtj���0� ֭��R�+�����������4]��RG^�����s|��U���'�W�������5mǞR]�`y�z�N6騚��k~�b�l�w��ΠF<�x��y���D��ͮN�9������e��5��l�7TQH��t��[��CK����Ax�ش!�a�A=>1����}'�h�ݨ��K� bL��sNVݮI����N�a�\;���uz�e���͢?w��1k��v�5"Ug�ZK�o��O�G�ud���\l\�kk�-�=ܱ�����hS���gq��l�Ї t����H�6��?�p���T���+ё�-�q������Сk��=y<������Vv�C��~��~��v��=��K�ń#�oT�)L0B��-�ᙯ��n�����w�z,2�l6�Ц�h$���^�Y��O�V�'�9��cUP�v_��18]����3�%}p���'�OtPYr��8�����2���>-�¾�~d��#���Q1+z���()Z����M5�v��w��mH��D"�ȩF�k���d.�/|�V�	B�1�t�xC�+ɤ�y�ج�����ʒ[f���{��͒t6Q/S/~��`|x��.�pV�{?�m�̄��$^'�C#��9��+�����w[Ǒ�U0tK���c��]&��"@��×�9������3b����@g/y�q	d:��������=��I������
T:�U�J����ޙd��p
�W��g�th����h�q�WTC��il�T�N�b�}���p�k�#խ�����D����M�jp������)�&b�/W�t�B�6@*�=����34\aF\����'cM=�Ps|U���B`�b9��:�[�N�!%��S��psd���D�4��tI�]L%�V�T
w�yC��U(W�?8I�p;T����-MI�G���<_��5�B�p�F1�t!1��Ś��	Gmj+\�S�������$E��C\������s��r��h{.��[J|���o���7%lNV�RZ��L�[�W�E.�IS�H�W�blܮ "l%��{]��w@����.h����N���h�L�﴾6YQ�4���~�w�`����L��a�)q�%��8��/[�a�4�Pض<cK���IzTZ�K|qU�kV��:������-#H�{�S��q�ω��$��&�m#�%����̈́�]v`�n=��-��o�f��� Cn襓	��4� Pf�s�Tmz��TY�DX���Ã}ڻ7����cu�{s�1�~�g'�"��z�t+����
V%U�+�ך�h�n���'�h�O�yh�oi�݌����bl��-9n���Xk@�i���� ��VJ7M��$j�r%�D���E�j�j���zJ�I�oU>��?�~r�d�2�ֻ��8���xl	�Φ��f��;Bx2����W���k�k��؁�5��ͫ�c>MJ������D��o�z�ۨ��1T��gf�2���g?7�I'B�cp���/t} �]��p �;8Ƃ���>�Щ+6�_��@0p�����Sf�b�&��q�>tMEt�s���͕��s�s�x�:M�(i��a5�}�i��}h9x�f+%Ƕ�f������hS��������������Mϭɒ�		o]� ֠69i�IB$p��$�ݒ�l!��#N��Y�)|����vq"�����n�a"S?�O~E���O�)��r?_�q�Ǥ	m$.�#��W�����5gh�Q�i�8H�d����$�>H|C�/=�@���������@o�r8���X�T>��L�!�/�KC�CU0Y�Q��v�jÈUU����8�AQ��1��%��q{���Ǝ�^����)fS`��mKъ�����
c��PR���m2p� �#���q���|�п�f�f��͎w,�d��|L�AJ91�l��|B���*(�a��?X���cm�:�Q�J��ԁ^�2�&}g�܊��CqAY�fã�O�E"r�썢�I$`�{��Elt�A+�vRW���\��o��I1�1.<��˗�b�w괃�7���	-[P�/����kfu����ǀZ�DΣ�u{�x�S[e��-��*��k_s��3�rj�-��(�7�A&W:h�7_�4��"���-_����/&5)�غ6;�F6�"1_y�6�r�ަ�����[^�X����A����®�(����� u;�ޅ�m��v�w�˾��Ç?�?e�����Y*a��W�nx��рy$&\�� �����������ұ�a��D�����W��|�$�(E�MD@F]�Έ��z��/ݑ�B*	7��-�{�c1#����/�
J�5�&�b��E�iiP0����Ꞃ'���=]S`�d/�dY�|5�:nEj��M���@`���%f���@�j[2��8`�=���\�슬_ɭ?�_ac�o�?d��R���$�O��7O�¥cF�i���H��#W�