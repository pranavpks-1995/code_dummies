ܢ{�w kb��:����D��
uPͩ����RY�\<�_�>���e����z
�8�  Urb����g��q*N��b20'Gb�	�98�R`�~(�9����c7iR���������^pU��Z�����&���5YIsUw��D8FKBb�����>��Tw����A��_!��
�'dZ�bZ���ǆcn�Xv�V�eIZ�jE �|���&<�*<"��o:�ޗ�7e�ir9��	�j����H��t�$��bE}#H��H�ֿJ>(ޙM-SP"��{�����+&gʥYʞ�K�p���ŧ+@� 7*c�Z��1�Ϝ���y-��U�`d�6�sIa�ٳ/������dCF&�(Y��5Ń{~�%�]���ǌ�6�M�	�M2���! ����PͲ��dKe���~�?�w��(R*�L�o��/>��B3I	E��*�M!�&�&Hc�r��c5߻d��Ji������W%�g��J�@r�@4�5�ޗ����ID�
w��d���_�o���j/j*
�VyEt�{".4$N4���t2��"��3M�����l���'©0X��^D�*�`��WS�Ɂ�f�o:s\�t�]l��W�Nj���9.SaN��@,���7�J�^b�A�O�Y%򃤐��R�4r�iZ��/du�s��kSmg���� 7����\�I0f?f��N�w%�~0~t���Л��?�`�;U��4�S�0��:|�n�{'���涠��S��N�兀�/�<5��Q�-��o�ޠ+$ٺ ʕ��!�Y^�=�b�jG��X�U���>�R���FCQ(�3%�Y��ϪK+t������%z�R�W|����jd��;_����d�IW��EV'+{��]�j{Թ��4��� ��������`-���H�dp��#��6�g#l ��L�&9L�R}C+Yy�`M��@NB0v��2��p��x�+]KEn��.��n/|�����:"GY�J�4t�'�/�o]�[���.�挮&�M|'�#5͹�ê-�޵�ϲu��18[��� N�?�L� 3��� �&bym/K�5�X-��,9���-U�/���rSմ�����{6���>P���o�AK�}>бQm�~(e�������K�r,k�����7��}:c>����<��RN���������EA*�����]�Q�+}%�-�ű.�;Õ ���&�l���b�Yg���#�ޣbv��>˿8�g「��<�X��N�ĂxJ���k+����йV�F�쐽k��I��:�WþO;�V8sD�`!$	��� ��0�㑾�BAC�1*cݤ�<�C�]�:(����J��Lz��5����\����`�TM�m7<�Z3�2�h���A�t��e �f�M �.���n?#z�͘�wu�����N��a�T���LV��~Ģ���>��c����K^� Z���0;*���B�`��_�}S�l!/>���}�ta~��Xf��Į4j`������âwQ��ZI��4�]lP~zЖ��8�#�9�����S��ʸh[�巀T)����L�RC�4��^�܀�w 9�e����qV#	F.�l܎h*�{+����)�Iul�pU�W�_�kjrQ�m��|���/(H^��A v`���Lsj�Z����q���/�jT {�އ�QU�<Ʀ�M���O%V\�)dwK�.�����3��I;�	��J�c/��7��#���;�T%!j{C�c�L�X>�K��ALҝK�!]�` ��+�8pb6�&Q��3�i�s\������4S����&�$f+�%+ιW1'׆Z����-�K�uU}��s2���nn��ܾ.��f�l�X�t��Jg�����4ձ���x�QV+*0{h�m�Ǚ �f�٢�;?=1�EKD:op�Ed��n�}~����JKz���+>�.�R4Y�H[���یi7(Y�ac��Z�'��tY���.��|v`i�~�*F��2�k���zNh+|t���d��o̙F�p7�q��jH�E��p5��ڴk��.vm�
3ΞpM�T��$�6'�)�����	����Ԅ'�t�e�}��d�'�O�x ����s���l�W��c��&��+�1�&�[��F�;��,�޹�h$ݩ�Cg��tz�L�P�j�!`�����=�g{�ZX��`��ʾ@<�[�����nh���V���֪�es�#Z��@��F3a)�M�K�Ik�W����q`H���B=R��q��������"|���П��N���id�ʰ:�A����}�mH���-ţf��+�)/s̻�¬�`�8��7Ͷ���ԸW����?����l�(YS��^5��`�W�����(z�K��w���E�;�|�0f����
�	�<']�`��Z-�zSy�=�z�~������^���,�#x��)h�u��>�!��R����ՙ���V��b�ԅVZ6jh��� �t�'�pZ\����4xFP�I51�H~��P.#���\#a2�zޜ20��`�$3_r���D5~��k�8E��hu&9��EO� ��������!��$. ���i��@4:��d�� \㭿���jp�K��
]��u��T�Z��
xqPb���n�m��^D��� �I��'�7�7�a�&��n�tH(��f��E*�>Q�KC�����
B�.h	�(��Dc��CKU$٩=�B���Ze���� !�P��� �Opk��Z���a�@�f�21��#;�� ��e�z�d�