n$UN���A�$  � �F���,t`�A��h"�`���x�����,�z{ Sz��,0����eІ����f��p#�GB����J�%~��H�d�ZuS��=`�[A(��d�`ĉ^���Жl�1���e���*7\k�����M����,�k�:�t?����6�B����k ۜ
����j]<��=�YQ����DV���Q��b���
�,C)��βd�GB3qE|�}1�c[�H7���V&zѯ\�i�˾��h��EhK �2)$�Y�����#X�OM�vޅ�р�\�*����)���_~����}s��a܁�c+>az@�>c�p��Z�Q��7[�S�9wZ���9��cr�!.�
CTf��tKG��Y͆���Ɋ��WV�XL�7���Ь�����w�.�f���}�䩀A-��D���!�|�������RQƳA���H��IC�8��[,-������Ø�\��n�a�)��f'�УB�w   � �-W���	�b�q$�!$���ZX����������}��a��hLλpC�K]ZN������.Z���}FvQ�o�7�d���K�����=EV��d����ZV�+	[���iF~��U������z̜R�kT�u����@"����sL�|��}�Xz�^ֳwt�r)Ds#͢�ѡ���RȲ��������!Q�G1<����q���s'��t����ʣ �E��$}�?
�,N�ֻ�����7���]��OǷ����������ĄȎ����!M�4f�Ϋ��d�U���Z�'n�}��F�䪷$�|wB݃PJ�i;��q����A'u��o�iNT5�i��p-���;#������O� g�~홸�&��~�J)++6��	�2�*O�X��Y�U�B��cF'�Κ��1�������H(-!��*�"��м��z^@�L�n�a�Lz�u������:�q��Ю�pN>�G�>B���Gޡ\֣�Mw�emp�EM����������!����!��Q��2ը \����yK �a	���u�e��=�L4ͧ|C�