O������i{�$`\'m� Y[ݚ��.��9��Ұ�9��Et��'����g���;v@U�@P�d��k�T�X�J\   �!����Dc��l�qUP�Ԃ�Բ �ڗ0�	�o���N���J�y�e0���F�,1`�ZP@�z]k����}UU���?6�ɉ�����[>]��j�R�T-q��T�ڰ_*s�_<i)^L:7��J�o�%��� ��v�EW:'� 1���!UM��G�`  !�����!H��a[�8e��Yu�  �\ߗ�+|����]�@ZP
F�ss.�2��N��Q��53$�-o����Qe�
�iSO�%�Q����Wބ���W��V�q�_?��XrqV���G6 ��?x��;ؔ�buO��u�2dt�q�o� J)��P	��5��ZC��d�@  �T!�B   �`�U_q:0Q4%L�h���G;�?p���e�}���H�ɮ.����0��U|x���88��*��f#s`
�q�����A4�P��ѐ�l�`�W�^���8ǻ.K�L����]#�2��U��sY}Ե�r�!׹�L.�i���ѢR��q�G:��Ԕå��հ&ɥ�}�m;��T�Av��TA�G�g�K�p�p,F�:�ʖw�J��l���I�a���m�'���̘sF�.^$��Y�����^�J�����*G��q��ۣ}l�nr��k��SR�A����^��!Ĉ�{��?2�Ti�4��d@r.�&<�鯃M��<�C��Zu����&G7���%Pf���gWJ��s�Rz�oGE6!��aRD���WR�8+��ٶ;aUs6%�9���5� ���{������ʏ��Sf�}����Y���!�Z4�$U�ߞvSB�(6���+^3�3�
a�Ȧ��c�'7����ro\t�6�6�_��չr�����)���t�a���A΀h4g	)	X�<[?�'��#`T�^����V����cn�O��-��[