�� ;�Q"�}۱�<��K��YkL}M�#��tX��-�w�y��q����G	lȭ�u��/�_�]{�aoـ��}���	,A��˱��V��0�\e��A�{�]�ڦ0=�ʢW��N���6R o���zdgs��ݠ�e��)��������#v�a�"5uwT-�ػ�Q�|�/��Z]�X�(U&��LV��
��⽨B�ۊKm�������/�5݆@4?���hhZA�y�\�w�GW�7Ò> ;����_f��d�L�).�_��&�lF�P������@��x4�G ���X����h�j�,�e�h�c�����~7=�J>�1���Uк3�&b�[@���b��	���Ա�퍥�N��S�Hu�B ;A�z� X�^Q�G�zFOh��qF���,��FA��
�ă�6�L�2��EC[���_BQ�"R��PY+�4^i�cR�GqS{K�S Z����/���G	�`8�d���I��5zW��#X��w��>P�u��#�:<�ֽ�(!�Δ�߮H5�B�/�Ȕ��F]�rCx������x���-����eP��⾮�)����3Q������Ϳ��F�����Geoϑ���y���mE&�r�A��@Kb�����8A�-p���`��Q,��՘�p�� [���8H�:S�#�(��ax�nk�<���=�҇{�ՋY���1[5t;��F�"�`�5��nhK��A��P��`��X��D
�La�&`ͫDyoH�G=g���hϥ�ŻEa.R۞���� ��ڥ��8�?�,�4�A��j{Äyf2&ț�!�~Z�Ox<�RΊ�%��t�$+pr�r�~fڽ��.�U�	�è���)���3P�т�1 �O��:�e�-�����c�w��d�M0�W���ܠ�
��!�ψ�t��eQ\���5�w���s��SZ������4��1.�}[ �yć�q�G�������kq<TY���@�������I<��������+�O�Y0�+ځ�Dkd��?ȑ��~�)ܠO������n�7�׌A�c
Sx�CZFO:�;��'|�Q��iف��9�:?�6Ĉ7ÃB�
��Q���Y���93&���<��\t�z���d��%|0��c�z����dB�
_d�R�3mw[#��S[+�|���A��L�l�Z�ꭩyGOG��-��*:�5��C�g����=��-�-
��ډ��H�{��O����\w-	(��H7����#�\��oH��:!$R�V�����/1���*���L�+*�:�H!�E��N���8��׹E;���p�n��G��a��b�Fy�eo�9��;�E�;V?�K������|�0��pT��؉?�-�oL��� �IR���73����v5Cn��!�t%M�pYS}	�n�J�{bX�s�B\��Q�M�W�@ok,���tY^K+�A>��Aoh�g`*�
�-��"����k���9�)����tZV�:|8T�� �⋫�s���1�rQ���KDPG�����~��)㙋���e���