4�b)�K��F�1�V�s*���ɇ0f;������oxl"\��nYO)�{EU��u=K���H�NPQ�qVڀ�����xJ~�-u��}9��~��������dΨ����,B2�7��ʟ�J<��#�r�eDyޠ�se&3�����N��6,�	�',֞4믔|t��[e�� �T������%�;ȫf��"���e���p�o�]k[�
&�rxg�����V�ב�����XR�(��gw�aT�u�(���Y����;j��kU�*����C����*LQz8&E��T�엷��5�G9����(l��У�j*X)���i�f�і���u9�(I����~ݥ�8V=0��/����<�� �����[r#�%u�|���/��� h
���������Z�i�2�,��e����y]�Kq��g�0�_�ҍ\��QԚw��F�ޓc�(QG�1Cߠ� ��=!>C�+-�mq��	�+��rU��$<��u�k��Q;[stk60�|�O&����Z�V�n����_����{d�LQ5�p�}3p��&��sC�/� ��fS�9��#Z��F^;Ħe$�CD��c�&f0d+��F���)F�+���U2w@��ir�<Hk���Bq7iM�|7y^���b��l3^�	�K���C�9sy�qCg����,�4�G{���$�W�?&�u��� �,[S���A*ysH��4ۊd�b[�s	���u���W.,�y��o���s�uCѤ[�?����,�3�l�9��32g򻂡(��-l��&�� P�Td����7V���2���/��)�#�����KӯT���|<�Y��ߓ<�XpQ��X�IioO�<hDO�U���[�$��ύ|���0�*��y���dZ��R��m��!�PHL嬉�<���,6}�mU�jt�Rw���W��*�0MK��~�+L�uނ�����2%=�y9�3o�G7��:%y��꦳�ȼ:�\f��<,����P=	�9���I��Gk+�/�=,m㌁�a�rFF��~�����<��E�De��%@����;��+�_�(�9XT��Omի.��HC�뵴�<�'��dU�t���^�BՈ�?N��ř���	QJ�~��j���|��!@1]��\*"w b�|�3�i�˓mPɛ���gO	�q#`�P���y^��"���<�����3�N�7|�~H	���&����
"��)R����|�.x�f�>yU���5x#�n"��fx�l�r�"G�r�S�=Y�sW�$>5,�s�+Y��]x x������~p5�@*i_O�m`>|'7��$��LqPVy|h�Ps��*#��z�n�f�u,9ƽkZ7=۶�����E�sKb"���D��TJ��Lv�L��N`F�y6�m�҄m՘���ު�h#-�N��T���j�hR�8�}�����v�k�0�G.x�P�o1=vS��󨡰������;٨��~Z�aJ��ˀ��SX(�DR�UL~<�;=�? ߔ��DY���\d��r ����͡�x�|̉'�A���<�*��;��	��
� >���S4I�x�R�W������@Y���{L<����w2$4��Hɘ�n�d��%(��&�Q�[ �g����/@�` $��)9��߶�q�+�_睮�a�T0�������U�20TH];e��P����FK/��!V@i���+6L��>dqsI��7o��O ��ֽ嶗���-�?c���%�?�9���}&-a��_��hJ[��eh�VѼf9K'Zx*�K�������鍫Gum�5Dp�ėm������M�9�[�fW#A<�k�`�� �̬kLm%}�����j߮x�`���Am�j̵-��0����x0z
̩��㉑?��δ�!�xE��B�t��\ym�c�WI۵]�:8I��EB��h�q����iF�D���=���Sg���w}(*o��=aG�k�}�;t��R�!S�ԳU�>�R#�#��͙���J��C�u�:�J�㦲����ȭ�x��)j��/q�y�� �'f�h