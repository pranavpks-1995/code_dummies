��f���"
�Ѵ	�*<d�נ�B܂ɵ�>_������@����#Gl*�?�� 3��|
����>�m��B�?��'��;\*�A>0����	�w�?z�����g�덃����:Ѭ5�l��+�䉎��L�mE�6��$�݇�x(xx*���a�0�.BF/	� �~&�(��b���C�#9�o��ښ[<�׸��a8?D�e����8[���e�򽨂!� 0���.�E���(�
�5d,i�X|C� F�T�-zXv�łݸ7B��
���ZI�!*N�\H	9$�T��_%�@���]>�a|llӅ)�!���xD��9�-������HlJʏ*٪���ID��=+g�/�SǳI]��h䩴u W���z���ax����B�`�p��b�k���	�M����q�^)
8 �uA4RE�;R��&"OW���da�L�7rV�7ı%t0�s�h��8���;�h�vJP���
�M����S/��`�s �t�	��ҳM	CS�x��4��)�eU��$R#�E[3����Kw�yd&��ӅW'��8�s�N�4�6f��{u��QQ�q]����Bfu�WO�:�Q�J6D)C����qr�f�^AZWj�L��zzL�!a1��G�JY��ޗDV��i��+���gɴT�ӁE
���p����̃T:O5�P���{��E�PZ��Nked�Kq�	�8kJ�,�rT-#�^V��R��p�X�(s	h��j�ne\��<LȌa����v-t^Ɏp�\�V�k��w�ʪ>���~�:
Sa�S�ԍV�LN��J"��~t۸u�u?��jW"b�W��F����[�O���B�.��{Û�7��fxI�����÷F�t��S6f̞���������