package generatePRN;
	module program (Empty);
	endmodule
endpackage