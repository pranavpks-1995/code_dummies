/?��iP����."u�7�%�h�
�Y@j��Ѭ�gZz�;nȎ�/$8�ˡd����G��V��3���A��s�������u2�7��$���L���Y%�h�?��H�L��;�����ú��su���c�&�+�َ���?�g���h�N��u,z���0�2���(�`{Q�ż��.���m6}j��tM���A�" ����BH��O��O���a8�v�B^J��ڣ���.��B��p��[�&���3ϔ�o\��2��w#��jG��޲�� �P��*��{_cE�%S'��]�ڪ�[�gb����̑=�ꀜ8n?[s7�%�7*�>��r�+�����w�qA|����>t�|O�P5�j��㸟��B] IM�x��w�|0�����fY��D�u�3��䩙�I,Ɩ��
��~A��Ӧ��&�u։��ʼ��S�ۧ�;:��rl%N�'���bRwq^$[x:�1���ݡ��0{��H����{�}gyTo@xnO$9�S��#�|4&��hr��ZF����h��H!�+9���P@Y��g2���{���Z~�m�j���y�����~PWfR��"�  �hx| �Y���o�_:���l)`�V^=q�	c��,�!Da$�iM���Tw;@&�1W�
9 �&򼭠����J�F��KM��9t�e�v�Y�R�1�j
���KH�<��)	l7��E���j#����tEB?�����Y)�����bٴ�Qg�|×B�Ts���ա���4B'�`� ���C�� ����kQE��#,�+�kP���8nN��eQ�rg����A���&N���kt��$�z���|4U��P�I�z��
�X�v$(<�Q�DHk'7&�S7sԣe����.`�;�b��淀�G�6��2h�ٴ�׃"1O�\�"u����]C��#��I�x_7�����Q`���?m�, ���$�h���Ҍ�y4=�i��R�	�󠭬х�@~#t�-�i��E�������:'L}\BϢ^Z��Z�˻A���(}q��$f���X�"í��n@��m3�W�s�Ȼ�릉� ��
�"�Ǚ�%ErYT�|��f�UNl�����K+0���N:S�;LTA���-_�C2���-rHn�ڨӰ�'�)AG�v��}���&�b��0�	bý��B�v�*w�օÿ,�g�1c�Q�.3:�Ь�<�D��ln�9�n����M?H��, �@���,TIiۆB����U�'��rA�8O�l#Q�`}��^uiyL�F���s>ԽW.�g�vD\��g�G~j��qw7��5~����?��܅���SG����>���4�S���w�x��^�y�(�zό'�e���l�����G�3�6@���E�_�r^6n����D�g*�.��u�3�Y��R՝��z�ڧ��Lɢ�\���� ,t0�]"�UyZy]8��6�^��%F3P�U�����e�18P��3O�����ܓ:��g��_�SԈW5����,��ȱ�}�j ��yS$�r`&��h��vH�ao+U��p�V���a}�R�6!��>W������dn&1���!NyБo���T^f���I��K鋌�.u�]AN�nu��T�U��M$����0T���*ϯ:��YC�%�G���c�/9���y$�SwVV�f��� wi�)�M1ţ)�4ХE^�+-/4Q���΃�K��
�#�xv@G�J���<;B�=3����K��[0�1gm��a��ζ���FE���i;¸�M�h���\R�0X�#E~���Ђh3 �oؔ��l'h	�[oA�W�h�#���u�|�۳`z�<a�z�F�EY�'E��@.8(��+���	-H/e��q���B~ͧ�;g)fiF��81ja��ͪ������}\m�Q^e��c���,����Ɍ�	�%R�:���ɷV� �Q�k𔹨�+�kR
Xk+� d�V��]�~�6�L�0���n�f=� _2$$cw�?
�E�g��s)�~B�C$$�ji�>��+��,*G�=��㌇2�(t��7p�!�E[~�a@��0���[��_Z�m�-^W��Ƥ�b*�*�L4a���']jXi�m�F�M��D�:�5^�P�4�s?}�Q�O'�@6J]
+��H��5�K+tq��T���g�v��DC�:�4N��q��2K� ��F%T>��U���]�IaX�Vjd�#�[u�0�r��G:܃u]����~S6�8�9L"����6�-����� �7��)S�p��O�Í�  	��%RW�c������f�b��s��c@-�P"�]Ť�}
�-�/��)f��ZX������M�ؔX��V��N@JQ����~G��O�/nݦS�Q'��b����5T�ϓ���|���մ������Oe\g�ۘv<ޝ a�^3�36"7��̟ک�x<�Hj"W���� �Z7����6��*y��\�b-XS�u�0%W��MgVSB�]S�ˣ�jլ�51�VHs7�%X���UL�K�l��DZ�HH�hOb�
�}l��aeh����4��_���}�7��t�t��*�Dw�7�v�U�cK���9.D�S(�DQwЏ�9 QZ����	/`*M�!=3������2�DO��H'LV1�融�e���D�Y�����+����"x�E���Z�#������7�P��d�F#��T��U9�cs�n]�&h̶(���bd^ɲ�x�.��Z}��t�o=�V�� �C��t���_]���'������?�)��M/��}�@�c>Yz�����#����%�b��=%m�{����j_�o��GF\z�Uq��]�8#��a�F�G�˛���ewG7�w�`hT�G١X�(� L��&��, ��T=\���z@ rc���HO�3���eAz�ar < �[!��SFQ�V�����wAS�����v~�:B_us��h/c}8 ������D�EH�#Zm�#�nbP��s�{~��h�\�Puy����VA{�ē�>6lz�7�z5��tb���K���5�(^j�k�(-%,a�[Ez��THP��l۴<3�O���G(���oh����F�GF��Pnփ���.Ȩ!c��!�U� �G�,��W?51: }6��j)j� �I�'
+P|���b��b��x����S��Bp���J�@�[���j�6YSM�a]�e�n�G&6�W�[�Q�:��@Ij�x> ӎ]��=��Ŵia&��6|�u�DE��ԙ�,�32s۔����َ2�\8/e2\��R��xVŬٓ*�FF�5iv�>�z�� wF�5���z�~y5]�K4�H�{#4 8�
���ҧ�Tf8��շ�ET@i���
�:T��*�f��(a+!��e��$��[�&ͳ�:\ߖ����BH'�f?�d�{g�a!@�����`rf�So��M�R�5��Ok��쿝;{%�7�l
%���B��@��?��r%0p���:l5���g�O��2/H��01F�'F��f�K����tN������CW���3��~�喟��(z����)f3����m�L��5�kĵ.~`�vEs"-?հ����C6;��T�k���ۦ�B��|��S��	��Z�d'.?O�N�LDN�p�,�uW�xq��H��>ư��h��ٖ�_�7�|
���bM\����xl�����fޠ`�Ob;��կ&Af����f�ٲ���
;I
-�X=��*�$��sX9C�~=
��M�$.�_��B�+0<:��*���.�Q�N�.��J���R4��r�	bmPP���'@T�M:y!�A�"��0d�����֫�66�w�Z��Q�j�C�O�pW$G���"g�dh�n�7_�>hZ� V����
�o�^;���6��@L1X�/f놯و��G�F�CFaC��D�k�����D3����s��\*��~�q�#l
yvt���h�y�蘕omue�4,���bĖ��k���s"�(��m(�oȧ�1�|��s	͚�g���[D=�����]����>�ɭ�$t����Nn6�.�jm���I-�5��%��L �
N)᝙����ӛ9=��s��<���Р��<Wo\wQ\��*��W��M��+0J�����w�&Try�q�LĄ�☑gq���4�Vhu�{��(�c$V�>�`�[Q�I.S2����ݼ�H�,�>_ �
�" ���xKuL7U��� ��lA.���wǬ�ς��GM贓�,4�RK�5�ǿ��V-�F�&�gEl#�u�6�Pw�u\>�c�� ���L	���`�G����N��p�a���&����;_�|x���z�T��v3iء�P8�^��� ��Ѝ#(���ިDJ ���E�\iǡ13�������u�آ�w�Rb��C����BM ^|���i�C���@m�� ��`7$�
��8��>��蚔�A�L��lc��U�J뜷S��t!�m~ ��$q������r~at|X�s.W�=���H	�c~�.Rڅ�}�����ZaJ@��M@ �ޙئ������|6�gM2�1�T�-��䜿���mr���!���輞��Λ";�O�{�7vy �1���R��N}�s�(�%��΀F����������2��x����`��(Î��眃�u��=����*�6'�5����S�L�s7�%��倔v�	��R)�����OF)a�)X{B�f���n�a*�0�IWI�(��E���  � �f���,t`����8�5�?��I��rG["b��k/��m&����^�
��H10s�C{�F��ٷ��[+�b�t��mIN	�N��Hu��1,FKW���6��l1s�O�$� (%au��u����M�ƈv���:�*1 qP��i2�^��Y���ws˗�Fx1H��\,���;e[E�c����1��W/Pr�%���N�Y���C�&Ub/�X3�8.y��2JR	��|���d�۠a/K���� �j��ˡj(�7�ͷ�D��'�S�Fh�����gp/�B
�F�gֈ�Y��:'4t�sB6%�2g+��n��˯s�g�!�O[;��1�	��Br!U�������)8��5��ԉ� �q�<fG�L ���u�(z���6����2������#:�F��4�<+l!� ��z�_3��Pf>������fe�o��ѩv�6�bĉ��~��yf����?W�LfH\on���Q'�o$y"�ϥ�m���[$�
���M��/o���C%��@��Z��Q���[)�ݤ2?��s���R��Q������45���x�`N:+����i���̀>;�Zǧ����(�8�'4��g�K����eS��CHJ��q�_΀,�`h��Т�Y��qʺ6s`���?fA�x����@5y�~�;��z��?X���DR�
,mN�Ў������w#�Ƴ�7� )O+�0��$#}�wǔ��q����D��cW��&��'����i�s���3h�J�JyO���� KL4��ݹ�fܼy�����{8bj�7i��u��_�ۜ�#�M=� � *]z�$;KԱ(��� a���]�kD��ġ`�#@����{���J��S�?��7Pyu��.�@���X�3����z>%p�#�#�g��x���4d��̟Y�`+���jK�X��$2ǽ�����Vٶ��/E*��w�'�l�Ď#�KL`R)��������ܽ�'�~����.k@��o��O�)�跥>r!`"F"m�,�cj����|h�@�I#Co��#�����bþ��OL~o(U!��zh�K",F��S�+��yp������G�����Ac��献[%���|ꙣ�*���"3o�,%��}�o�N�Pd*>WP6#z���uR�#&�y+~�+�lE���}�e0H��{zm��ǭ��~�S#o���Cj����\;}i`"=R/T��p�MR��㓕����y=0IZM�?"L��E臭�S�0�[�2+Aj�S&���%�\�*Y�adtt33L쏲���\�z#��\hLE�B;�ڛ�ռ��m��6�1�Ze���Q|�>�cW� >�/�ؒ��n���W��V�IqV�E�=n�R﫜����M��q�"���5d2���0�ٛ��JG[WؤأF#�"    �-W���#Ѡ�b!C^���Ŝd��ABx�܎�G�ٶNvR�8�8<��-�fx��q��D�=�����24P9���E�;Hq��z/.!F��iy�,�������2x&_�y
`R��2� |bS�S:�a���̓c]T����0s�.ȁ�0���v���[�r'�uP����H��\�R�!����ʨ6�i�9�2�76p�zi�|���C��d>�h�!��Q�:�����vՀ$�,���}�
�uϟ(�<�4Y���vd�}�B|����b��%L� _�����K�
ۧ�2�d�{� �=�g2��Bjs��q�LSg����v!��L�J�mxX ��X巠�Do���as�	_� �Θ'���jH�$���|��H�3�9��v�n���:�@K|�Aw�2�,4h�V�KSAĞJvRsb'�?��z2���I:�{+�����ϝ����4ǣN=��ĎM��]<`f�1��5{ގ�#j2�u�B���'2x�TH��C����r �J��x.e�{�����a_�t��s}z�Af�K�Ͽ��9i1��^5�\�������6�����e�w���^4�
tF��P�DAػӞ�1��t�U�3�/�g[`��Y�l��"�.��B��v19���}����Y�� ��X�Y� >����WKj ���M�X.[8���p��%����ԥ*�f���Sϝ��<���Z��wT�p%S�g���N�7�U��,m:^m4�)*^}��nt=�0P��hYjI�cQ�xbj�y�?�\�+/OM!_4#;�0F���}����g��QR�,�^z��h��F�Pd�^��@�<�It����^x�����fT���^1T�z��=
��d�`.�)"�<�X$|9�n��~�!4�rF���1H�s;<�FH�F�����d|�o�r��Z�u#?�]��o��q����إu��پKTspy�j���3�ڳ�Ky4�cΗn�e���|�]m����!��˶c�vׂ��^���*�D�q��ju�AK�o�:�O�C*i�*��9��K7\�J�,.�y㚎����Џb� Es����1�}L:x��0��-��k$�z4,G0x�����J�*��D���