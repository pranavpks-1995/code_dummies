�>�&�	��}�����]�A�>T���̮@�� �i�E�q��{���k^m�X�e�!�;�b��F��ˁ�3Qݑ�O�k~E�6�q���m��ӽCY��e�l���[�hޛ�������.g����!4��4<�`�3*8Y�K��F%����߶/�9@�g�����E ����Rj�� J%�=:�T?/�B���@�M�|�?�0&�E�e�J�G]�*���d��a�JF5��Q�#�65�=x�H(m{�E&�'�j�����|�� DV��n7��e��O�mE���y��]��Y����9>]SZ�gOa�n��p�fZ��(Z���������(p�#6��B`�FQe�0f�������+L�'�baC��ط{�l���5¡1�ݜ�W���y��,�KE��*�i-�j�=�����diǒ��Zs���g�u�X�� i��v�Q�Σa:�":Ͱ��߆�,O�����W�Kol��JBwjQfп��n�����,cd�"�-���$�Q·���4��p/�ޫ�4�_�	�����!l�'K@a���8�=ϫ�8~��1���N�EE��gn�7~C�jycW>��f�7����u�j_�`3�n!4*�يi4ڌ��ۓ�� ��C�܁�-���y�f��R��*D	��&�p�X�#����Ě<�9Rӟ��!�h��rdi�٤�n8BIw���R�J���3�)��oT�����*U��d��CQ�͛(J�