r��dt���X�B���W
o`aA�C0W�W�|��o�����0�i-�$�+��	�y��8��1��idr�5l����F�:qFj�Kj�W����fh�����'4���
�;�UND)��_?��K�"N������as��n�~
H-Z1����g�|�M$��K�9�G�}�c]x@�i9���H�f?{�5�*ǀ��ט��j���Ae`L������j#���}M:���L#S܁����ӱ��4Q6���v�Qz��%��NB�Ԫ�Z�B����hfL��+��j1�:6��#�w���OēA��#����=���� ��Z��Q}����iK������Y��?�<4�|[�(|Sy�S>�텬���)�&T����4�zvS~R5p����/����Q3�# B[&?���'x��H�p!���*�l� ��!QM-����wvM_/7�`�V��Э���-����3�w�� ����p����!f:�����(k�,Ȝ��֎�";˞�&}%�!,�� ��+�3[���׫{j������mZ'V.i-�j�
T��ϙI�i�V��a4���o�����.�ϓ$��}U��
bL�8��P�����ҷ�O38��Ξ;�pފe�br����V!�;ȜN�w2 �V���
��3炿�3G����Y���K@R��<2��	�L_m9�;f�iʘ_���m�ad�]���P?���V2����AExn?[�q'���W��*`�T��`�孃�)��X�@<)���汢�V�u�3�R]R��a�S��ì��gf����o��/�V1�k�@��޼@y33UR�^����	n�k�:8�	֙�Y��N����������ؓ�����b���Љu��� a��ĦC(����8�KQ1�$1��;mY��	���*s")���!�P̗�^[�����1fX��A�ҡ�ƣ{l�q��\'�`_�j�[%\gk"Q���=]��K��B�,%�S%�\st���#�P�dU�%)��M�K��T XU�"|u��I��U6�����̸�������L48$�Y��a����?��W�CX�����z��eQ9c[-�t�rI�}�"�#������
bL/����a����e8H�h!K��U�IٓX��U��-����m}e@p�+.����A������ۺC�Z��L+3'�Q�Wʡ��`�JA����e;
�#�X�c������^�+�EI����
@!�.��[Fd����V݇8�I6U����ܱ�󇱂(#1���Z�-/�?��S�Q�����?.�"�z\��?S��S{��h���bs�zQ����Ԫw\�*�v�`���f\x]��7�7u��D�U�?aZ��i����kJ�Z��J�i�{�.'�3g��U]O'����?�b��������h��<���t������'��K�^�J�c�mO��^�ZՇ�\6>n��iK^�*���\3�U�S��|�bU��F�DmA�?����{��-�� ��_L�sR�=��Z�v���6�Vr��D�Ae�D	�$    ��-��c�''��Y����:�@�{�����7Uۆ���������e��s �[���c����԰����S͛��e�%���x�)!΁ĭ�&�W�dF@ ٤����^D_D`j��l�?��
P���D|����z[���I5v �$灲�OL�Q6����Ӫ��u3�	`��L�������>v�]��HMMk��~T��.F�Ы�"S���𝛢_0fzi�W*X�b�.����P�w����v���:��W�'OP�xX�f����� p�(-5|s_�M%�ג�P�31o��xZ��Jq|D���L|Nt˟8e 6���6�7���Ya,c7\��E�aж>n܊:Yȭ}z�e����̊]F&�s��oD1;e�~�ُy�8�gdH�$���*�J3<n[B�s�*� '��q}��	�Z���֜�>C��2�z��Bջ{�+%��>3o+��9D�ܹ!f�M썢���+��NS}ʇ�UU����S4~���G�?�I�_/����o�>k ��_x�Bj��C��V�-�����NR��5\�G��&���S��J$&X��B�O$[��s��?�>�.����y3���	Y8Ş�^n��d(ʛ�p�?r%�n��$��@�d���T'���9�d��'����N�֧�`C:5wO�<���ô'1sI��**��	�r��"L�ݙ��h>��J@I�G!j؎�F4��	�lB�k��z�b�{#��B6f6�6����I~cM��&�aZ{�K�=� Mn�ȇ%��30����
�[�ކh���M[&7��q�>2F����NEFħ���d\�g�����&>�¾�]�\���� �~	��:S����s�	�	]�-�ې��=��r�	���1]R���ә�L��h���ێ�|���;0�]�
��e�Ϯ�y��v�Z>���.�O'Z�d���2��z�G���}�Jɼ�쵄�7fo����v<~�A>b\6,��-�Ӵ����cZ��g���x!`�E\�c��������!K�M�>��bYcHJsK�
`ށ��{E���ׂz�(�N=˼���Gm�ϡ�ns����Ӎ�t���5]�
-�a6
�ƒZE�^ށdx��y ��.q�����E���� �s@�G-	�|��f��L[ [�$Mc�vD��Q8�{X��R�ڏ_t�xD;"����zB�RV�   !y��@T�`��+� U�q�:b�`:����Yl��$�)F^8wlQ�����i(��Ѥ����r��H��H�Dr�.��p˃���ȴ�Cw3�zo���A���V�PE�1Q���r;Β� K� ���:I���W�I���%Wr\���чۙ� `    �!��
��Xd�P�Ul@�@28V����H��v΀����/eǈ�;<e��[��X��O�͏�ں���=y8������v��un4�c�h�~A��OA��_����h���4�`��,
��4��U�@&�� Fыx>�c7U{K��~�jWS��0    !�	�����FD(�XL�)V�k���O���n��ޣ�SX��߳�;Yx\q����n�R(((DD&�(F�12�&�"$�ᔃ9��C�2�݅*��WJ`Ղ\,;3�J�Y�x麶#���  OlDI%�&�3h�E+C9+s�Ff�����@�{|��	x�� |�`�'�۴�;:�7Ø�  �8!�Į���L�3���F�Y��׿5~�<R�m�V�3uTR�
9�VJ +��`����r�t�d�r������>@7�9�ZW�.<��!?���=�@z�x�����z�$��|ۅ#���c�TЌ>@ �'H�U;k����-������ �   �!�̮¢���2K�, �6(  ћ���Cg*3�W��yWH�eQ�!ڒ����� �ޠX( ��8@+�)�V�������p��ߦ� ��s@� � �3`kzW�l䡗A��>`#��U� n��0Yd �YB
�47��f[��~��ڀ�  p!��GB�@D6La��!��QD�U��GA�I���thp�?���CW����+K��kp�q�(�7[������`�#{���;�U|:�rcq��b$cQo������*�O&�N��q^4�
��6h?��d��P����϶t�#�V�}�C�l36w?\�   !��$���.{	%a�&��Eծ���cG�4�p>D��T!3����pY=�|n��`kq�;�{|�ND�6���/C���!f繠"j��/:��i���  O���u�^�]�  ��.,PPf��^�V���`ۤ:�m��f�� ��W��   ��h���q:0Q���V�U��S+j>����*�}q����/�����c&@�����.T�s�5H�8�z�QWd���tXUYf�J���DQ�sx��ڦ�.�����f�#�:��@�Τ�.�TX".�w�LRϬ�!�))��vJ9̓#�ܴ{J,�m�j�	e�-�r���ejH�8���"�q{��`�.����<J�|�`�r��c�3{e7R�Z�tD��Z��X杢w%o#;��\��ؒ��|%���ȶ�tH�糆���ȳ���I�����j&Z�:3y�0,VCg-�ܸ22=։t�7㋱�� ��4���W�X��w�����Ӣ8%�B�g��>�C�\��\�A@�.{��/
�_��G)��*���5zP�V_������]9}��{Nd�CKG��<����N����c��n����6��^�b���8Gy벺�\&[�^X�j6r^$��`}�d*�k�zE���gp8�x�d�"���5�'����[J�u�I"1.u}��Ca��C��[����Y��A�	��(˶�ݦ�?ҐE��c�5 �@Og�X�ݧ���`�N��)頡@	Y$ j����\>i*h��u�</ �#O�>��q#��&��.ŕe�-�p�k�v��ƾ��-���اhf��$K�ӠW�V�3��Drv�v����,�7�=�]�I���)�H5���b�%�[�>����W��4���4�s��60��\�]�t-
�>G��?����2�Pz�|v1�$�{��� 6.��K��"�}�w��LtL�~W���	៉t&r�`��-�K�������O��V���7�̓�p9�����ɨ~����˲ςI���%����ʈ�<��2�chb�2	�F�^�4 U~rMi؄���(8���T�9�?�,Qn8���[5C������c� {��c�c�%b��gqS[Ve� ��\����#8*��:�	���oN1�Mt����:]��F�@���/�����R��'X����_��-����ht�;�c�v���l��Y�6�J����e�黍{�H�rZ�>�k��{�C0St?�/W(:��<�LԘ��tT����j��p�p��c��*�����'��>�}�qi�������VL�\���{yFr��8�Y^���lg�L�X�!4�<��d�:]y�w��_��2k��+W��>'ţy�NN1w��FGַ*�WKK�K�5瞮�d-�Kƹ�	R���{�!���)�ıxg�hݯ��|���!��?�����^�S��UD�E4h]�l�Poի��D�t����A�V��8L� ���g���DCg���|����D�bθ�ר�uw19��]�Z��-w|��~�������`�7o����f���$�_|f�{���mN?�?U��
V�����ͩ�����)��v�F��̯�7SQr���{���f�H��@�]����KF[��_mre%�R�t2�H�i>�1�[�Y���һ��,_FHJ��i��
'�	
�O}���J�,�����K�E��D6��:+����c�h��~gT-%9thV��O��
�l�ګ�l�cy`�L�S���6S��H���	ۨ��c�T��qB�v&i���tg��&�H���tDOI{kx�i��|H�w�D~��wA�0��O�&f�$�#�Hg����4����Ū ��+��>'"�W�<�A6Y �5���7RW��i$���)e�¿#�sq	%���P�)�i{��s.��J��q#�ň��B���QYq��T[�?x�VK�N���m�8�