-
ғ��]�((/2�t�ö���O�����ܯ�6����
��_5��܌� s{��>F�?�?�k�6oCy����o#X3�k_�Q��D%1��|�+�����/q�l���p�ty��O�J�0�+<T���]/�|k�挣Y���F�3t��R�A*��'<����� �ҭL�O3L���ïC����.٪�x�[�����)�g�"��^\R ��,�&T[1+m��@�T1�j-��v%�i=�u+)_�c���&�*2)fv�$� }.��qu�j�D��RK����m8�#�I#�ZP�UG���;�;��.���"�X�JZ���c�9O0,�"���~c&#�T�?xȞ��A���`��������IKK����T%KNo<����Y+ _�*��Mmw�x��׈���<�#�[@
�vw�4�;G�m����gq\5�0��p���%<�fn=���1� �Z�'r\�[ߢM�k�(Y�ª�e�s��ga���˹Y����^�!u�Gű DJ��~�@K�Sv ��Hx�~��R.�j������t�R0q��@�:v7�t2�l��\̫12����������r�w~4LD��f�1"���έ�N ؘ�����ڤ�����$)�=�ƅbG/\y�S�um'��P�HG�0�� �n�O����%�x��1Q���.�T�m��c�3����(RK�6�(���G���=ܹ�?�v�C����s%t���H,&'"�u��o���]�r�XH�����-��Q߸�K%s�$���'�t�HTyH%�<�B�y}�ϻ��ҍ�Tl�|�0oj]jS�U�C��\ǳ���P3�Z"SU�B��8�t�>�~�t֔YS;D��/%���́y��7Q�YY�����Dr;-z�\�֗nTt+�B�q;�}d����n��~�R~\�k��İ�W�_0`L�+�V(\��j����j8a�����g� =O��DQ�����	)�����q?�R n�`N��+��t��h��n�j./�5�?�?�H.~��o��W�E�0�h�q��z��u5��B�ǥ<0�DW �o��hg�o�H��kJo���qV���Ӱ���9����n ߧ�i���,�YJ��n<#��%��_e,Z�$6�'浟6��ɈՓ��wK�h]�d��4�s>.V��pM��,�
�g�D'�̴ ���Qv
�C��08Y��O�����ܐ���j:����0����/���E�P�8�C�z:u"�y��\{�֪8��Jx̊8�&�P|5�B�R܅��j���-,���PҸ�&�I&��đ��Biߡ��V��`]b���eߨ�����������i��9�EqJ��uo���;MQ�D$�����J �W�_��7�%"���ۑZJ{�7�C$}���0x� m�G��j�+���������Q���Z� �2�1�#��u�ݯa	| �:��9�O8{��#��vx���ggmaL��8�.�R�Cf� �s�v�j�_#�^���QeV����k��/�.�rs2nX�}� �Vw��#V
���|��cJ�ǩ6̐��8l��((��� 0d���[-���nm|]T��-T=M���X�䩘����>⑍�㒜13���D%P��=����*d����-y�V�-�6Gg�wK���V��Nݤ��N\M�D��K�8�@�X �6O�x6�9dp�2������	�i�~���hT�q�L�[�>\��^(��ZČ����S��*��1'M�e?7glp�Ϊ�j�Z��t8��|4R.)���k���"U�h�@�)�إ��4����-Cܦ!�ڧ^t�K�C��<�D`s=��N�ꐵ�]�%Y���J��z�D��n�|�Mj\y�W����z&9�D�+O�쿑D�����G`]�ـ�?�FUK'���2���q���rܯ�~ʙ��EJ�s>��j����;A���E����m�*Y��sx��+σ���^,�	�|��UHާd�^�#��og@��)��h�7��N��*�V�?|�h&��b���=���%�� �����U�-$���U��r;��,3nΑ|o�/E���/��Q�>}VB����,g�zA=>�x�*�	XL.kV�rYJ~~;C��N'''/t����9C/ ��K�u�d�f�$b��$��|������G��w�8�G9響)�V��jd9D/����۳M�+����D0��G_�$��7ofwI![�rJֿݎ�ɩ�����/��k��Vx��L�"^f2L�O�t[c��%e�+;��rx�?@< 0���D�ڗƆ�"�v��j:�HŘ0��0���������I��j���Z��|VSIش�M�8�
˝�>�'�Er+���Ȣ�0K�گ��^H����<��a��ȷF��:qUf��x�5�uճ�rp�L5�Ć6 �?&M~���"����B��/i��-p�\��a���[r�F���u� �����McPr܏(E� �s��O8�&���}?#��P>�7�0duȯ牚в�e|���"�e�Ն��'SdÀ�F�4#�5-g�B=U�9�_�O�d�<n��fMJ4���ϏI8���$�d��f�FV:��$�l̾>�L}[w�[��c�4�se�O�p� M&s�i8��x7���r�ܴL��9�mz��'��-�88ݶ�Ġ�ZĹ ���� �b�V��Ool��aĵ K������
����̎[�Kܠq�
l u^�M����K`W��ߐ>��X�N��ۡ!=�O���}mt�	�+�	���m=���Gl���ѵW"�g�D�9� ��������:xNq�5z�э-�������مWw��h�G�Fspڒ�E�!�_?}qQ��1�0�X�F�}���վ�85z���j������:��)Qb-I�#5T�{l}��?��MGD�H��e����e7�����ͱU��"T(_>���:/����NZ���N��4&�Gnk ,�e�#�R��M܀�bR}�R�O��ɘ.\ྯ�ۨ����[z��'���r�崂���w����\�AP�%h���W���W�s�.║�{I�N��׻�9|�dץ�W��$�d���(�W��g�"��Vi%�a܄#����J{S�� ������	{-�
����U�ux.U���rX�ĤOyr��uM����AٿC���	%R_����@�����0ʅb?���sP44�����5�*#j��JpA&�X%����Bg�s��FYs�Rr�ť�}�l�qY����B�D�#H��H��%i��Eӎ��WEF���Y�㸼yc��⽦�Ѽ�ݼ]�(�ܐ�}in�%u(�*��z����=H��lH�̃