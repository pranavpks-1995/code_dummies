%�"ȱ#��kL�i=ٷ`=���l��@�6i�����acx�����i�u̩a���p�-F��fJ^3 \L!��������5���1�v�R����$��x�I�J�X��FQG��H��:q�V>��k@�e�X�]c��}�kR�a
�A�w�n�&��j��>U�k�;�����n/�I�Ԟ+����{9�$�g2�}<�Ԥ���7��9(eӪL�ќ}ēUf5p�m��A7D��Q���|�T�h��Qcn�+$c$�B�����
u,����6��J_�aI �G����L�њ9f��X�^�ώ�~O�a�Y2�%��M�F�^[���(�/yq��@��(�; �XCbl�tsژ���M�q���Άm���ǐ��'.I��KQ9@Af�-��� MS��Z�S`�(Jm�����x,�|�҅9����Q{g�JB+Bln��>����u_��,{��)h�;�����I�[�c��b���gM�I�ݱ����'��`m��=�e�klΰᔷoRˀP�R�ы�Y���yk�W�@�6�Ӭ��J�?��>�2����� z�@��FC7:y(��{&�f� �"��30�i�?���-�\�	ȅ�̳�u��c�pl/;��=�K�-t�\%��[��i��wf�_�W(a�=�l���]�$s���K����7�_�Ud�B���<@>�<|S02��aBO!���a^ʲ��.��2��x?t�~w�C�?Bˮ��:������A�����Q!��T�ۖ215�LFX�+;�+�߻��;�=6�A_��.0�OA���S�L9�(�=<nId%��/���R����W���nl$`�A1ꀒ������w�e���iS��_�@/9]&��V��b~^A(QƬ,�)	��wi���('��������%e��ؗ��O��ԀΜ��Эr?�@C��x�Q�O{}�`����Y/���+{awZ�dg*_�l��W���B!�{E��j���Y�nH�в����U�j{e�� ��G�J��7���%��Y
ġ=s�f_��LU�����j*^��ƿ��N�E��x��~��Ǽ/�58@,&s�'��<_����5���S�ϐ�_u�	��F���ZpN=�U?ڗ#6��&6h������v�ޮ�N�\Vbq�w�L"A���,(ޚ��5�櫍��P�,T�C��}�ii��\�w��}�sޟJ��-����1ɩ��T�(j�ё�#����g[W�+�:���.�X�U��كA�s$�qЃ(8���*��
���b�Ν���+�}��z�y�ۃ�,?�wֵ�����X���(��	�������@�����~������Ð����id���_XF���; �$3!dݠ�^�I��O�����2��^x�m�(F�2Z"���`��/�� �.<�x�Hnky���}΅p�($�
�ق0D�e2cy�^=��E:nѾt]�U�e��t]B����>J��*�� ���3ݔ��_���}.���$6�n�"�ݯ�H	s`m����cy٠m�x��H,�w�B�ꐺ�#��c�U
s+v��!�I��.���\�=v@m��w͵�|�	�|O��ڜ�}�1F�����D�>�LZg��'��&��!11�³_̕��#߬Y��z&]�J3�C�I`�s���uj�ף��5[�?s�n�]F��e�^?���RA"�����A�b����0�Z�y��Nԛ;{G}�x���dlL�-ҋ�u��}L���𠪓ԑx�.mG����y^�G��_���h�GC1a%�y\��D��>'�i.0�^����� \�A��?�j`5�EGp�iڷ�F��(q�G9Z���m	�!�?�����'M�<�Jl;vA�L�G�6_�"���KS�����n��a�e��Y"����;j�rw�T&୐��s�1[�;��>5#B~{�U�_0٥��c�3�̺W�l����>�F ��r"�,I�P�<x�-sT����@�ƙk�%��� ��~ul
m��ސ��yy� ��'���0^�O��r<
!sá����Y~Z�~5��D�m�.cuбi$��3Z�klK������WCH���v'�j�c/�?�"�Jܴ��*yKJ�V�v��'ˆ�s� w����j���ߣ�t"tف	feЎ~�qPgxu߃M�5�\�N�/?
�9�U��yI:��Ͳ�E��������h�5͗����!�N��n%,�?�8h��o����k�I����%oj��cZc��G�]��� �\���"r6^A�߷9C����ʐ~�B��	��..:���Sm(�� ��N�g!1�'�صZ\ă��M����y���g1�89z2�\]m�S��sH�ѿ�:���6�?8���?P�d��!��ϡHـ��WfɊ{�t�p6�b��L��ZVL5w?	�x��y�ث�.?���VX������ �U�z"*^�Q�K�2�m�j=��o���:��=T�R���1<0��C٩����}����ʡC,�r&�6��C��F�@��]��\Ձrݛ&I.1:�/�!�M���V��9i�}9��9t",���U	>G�/p��:�uQ��̽D0 ؗn��N��$  ���%W_q��>�d��� �.;�P4В�<w�5������/FR��P�l�x�W;]	 K��<Ge!�\P 8&�,�y݄�@�~��r�e_撓�XR2�'����wj��*,�3@��1�?��AI�j�BjA��Kajd�����잗J|�Â�A�}�혁�& |7� <�+�M�"5��r��^ �pD����5:��%�'��F,�?0��D��֌��n��7�`nNk�Kp��U�'��k��)��C�D�h��'t}=��=�ޏ�A�՗XB��>Z	`ĸ�+2�@jc�L�.!t�t�I}6��m�-}j	������M����x:i��af&k������^�G~�Ox}dT�_����ޓt�g�n��Vl��j�Tʍ�ͨ[��UX��o�R��0�QDG5�9vw��Rr��]��ٮ�~�Cbx"�ķ��gM��0���W�Z�� �إWJX�E��<�2�(z6͡��	����0�����$��L�IV�'	}Vk5��l� 
v�N���*�JJf�مi5�b^�S���1��dV���o�n"ꎃȺ�,NE��0q)��z�L�+�d)jl�t�E�n@��^��ԡ-�fL�(��~>�oZ/�\.���.��>=����R���h�L��Z�ͪTalx��S����bZ������SªI��#��/>[F�9�-K1Y%_B��]��$F��0ԺO7�%���?�|rX�����iloe���Vt�7|���/�$��s��4������۬XqSіB��V��B|^A TG��j�<N �m恶 .Xa�TeP��֩�=�'TgD�ޞ2�(w�N��E�1�I���*�m���Z��ۉ��G��ύ�Nu�z�C�%��M������.)�o+WnT#46h>�3�QDu���S�Ρ�ڤ�CP��KE��N������*1�m���ѧ#WXϠRNڿ�g�O�{��B9_�_'s+�₋Dz�a��X� .S�]	[q�&q��ssH�~C"(zء-���m�E���1[�&_���;m-�$)T��G<L���c"�� ���0�@��^{���e@h����ed�ϟƣA+���Ӝ�񥧌Ǌ�y����D�c���F������Ռ�J�RN2�s�����7�^����7��q��_j����m���$V�]`!�x�f���Xv;&�Bs��W�*�L�q3Sq8xm��ț7�Z��ߏ-�A��p��q��~�@C�e���_{p�*���p�8���f�>N)�����$]yx0��v$�B�D(�.��S�&�#i� M��l�j���-��-�0}Ջ/`.�.	��<��d��\�j��{�@�����g6�^p���N'0[��|�ڳ&\���묆�q�*���kь3d �.�n6�J�=`�M�����\j:|���N���4z5���se�;�%�8T�vR���4��bm<0����%<�$@,�c�:ű�Z��L�fIa�K�8��2��R�}���0tX���H��t��!e��?��v{,GG���ѣe�M�5L����hW�d�x�d,R�� �Cy��S{��?5O���{a�p/j4��t�*"� �ί���8T����ID!o����V5M���Rk�~�o&��YYs�\qn��Wt�4땳�@�E��%�\���x�
��Jߊ֗\��o���-W�x&!�,i��M�5�GX��<�ںL3R�������񞱥��
�^τd���I����w8_��,9�b�s�Gdy_���;Ԟ�����JbI�� �F�F:��h�1�qY�Dm��S�c�4�`j��R�i �w�Z@�]oX�"�Gs�1u�?��[�o�C���=�c��r���P�����6�%�3Hsّ\ۇ��Ņ�A)����S!�©���$1�y�u�r�Gz���Y�W# �z����a�z���q�p<2ͅT�H�����]��τb���Ζ�|�?�����`���*����z�T��K��-4m��p��l���b6M����h���1y+�]��3�F= b�3I!K�ɛzu3_ּ�vf)L{&
�)|Y���_%)���b�@}2GYF{QN:G�
cA��-'3j���n�b��<U8���;�0��[���Ӄ���L��6�7�m�@6sF�J/���DF&�2/�N0�k��je��TJ�j��M�\#dc@=���A�֒`�
���\�dX�vxu�E�-��ȓ�DB�ln�7%������5K�DM��\�|nlz�n�C��OUb-o�8��U����~��'36;Z���o�	k��i��,�	���:Q�J�*��Q��p�ܗX�}��I`�NH�i��)�S|�*7&#0y�������.1�/���)6�	��5`/\�[��R��Rc�J<��Ye#9	��Vc}�	h�.ĭ�h	�����<�i��Dl��ݠ��g��ֹ�'����Lr���eB*�L,��m���[u�ρ�p��#�a���Dh������_�,����%a5�dݍ�{im+ԛ����>P����w��[I�ٌGF_�:֙��<�7.A?����z�]��9<�Q���Ihtrc��W�}��V{�FQ�"Κ�3%�s��p6o!{FH�A0v�o�<�H�wa��u;I����!����t6�0{ٛ��Ư-���}k�݃C�KTC���u�XrV���Vv2Ε�1Z˓��cd�̬�M���7�*̗�Əӗ�M��(�f�3,º� �n�6��?�I��ԓ���
����p���E�MS8�=
h[�\)ˉTb5vw�5���%C�t�]&g�$<(���%�TAPW�H�&���^]?����_��њ)���|��b����)GMs���4t� He8q�	���y���P�c��p�M<WkP/��%�i
�����FEN�5��Zզ�O&�1S�s��'"p��]K/t��?�� ٌ����~�B�1���S�aƭ�3՗���H.&�A�tc�U�`��ǅ����42.WL���Q�L�BA��U~���'~|�Y�F ��ٵ��Tޑ���05�z�Е).�2�!�	)��#([�bj�)�1zB&�Yr�)�h�0Y���'S��e#ME��9��P�G����#S�#���<�,ʯ?|�=�]w�5��[Z�o/@جyj�����v�|D�9�:���?�K[d �x��6��,����g�a�g�Q��hl��eZ􁹊��_=j=z����y�eG��F�����@���o�N�h�5cl���MO4V0 ��m��BS���7�-a,��p�g�xd�j_�a�ݫ@�ik�?SQ6b{Q�����x;�6���%:��>����d�>��v	͵ݳ��[�w�gE�8lΣڦԲv-y�hw� .�"U�Z��C���iN�*������>haw�nq�� ����TQQ�XaZW<cﹳ,<�\8䭞�1)[dK��� P\/�����s�Te-������n�oˆڣ��R[�^8C��Ƙ�\���"k��{N���ͼ��sS�D�+sZ�M,@���u���Rk������{��0�Z-Pp�j,4��;QX�*�)Rq*7HL,�3ӗ�������S�%�T����[v4��
0��Fin���
^��?Ȩ�c)��V@-�;���]������&R�;		=@,�X�S3F..��r�갣H� �   �����,t`���4MG��W��G�(�D�l�ߟR���~����� {��njfI�%�R���\a���l-4�P3Y,ƣV�!�Z��5�#��lMUq��aQ���Q˭��7���2���+��#efH����z6�s�[]6��x �S��O�T[+��S�s�h�q� _2&����1qk/Ŏ��x���cN�~o7F�ޮ;���R�[u�p8e\��v��c��x)]%]�? a�������7����~�j��M�6�Y ��l��E@H�����d,�3������01�N�;�*��-�	4�֦�d�C�*^ }\G�n�k��U_&���=�#>i8��i|���!��l��F��U3�jQ�&�����i��F��Sr��b��ŊO3�'��6�[χ�W��	����͎A��*�A#�<�b��9z���A��������������z~7{��]�/�9-��羑Sa�@.q�+!��Y�K]�y��;��!���br-ã�����/y����ZA.3̊!o���{g��X���(|�����_6<� ��tq9�x�}FX\I���<��C�����u�z���B��M��5x%c
�d�� ����.{뀆"��|Ւ��@��XG˩ܣ۪F鮘x�����ӡn�ŋaD[`I'L�`���_�L�L�ݏ9�n��6����.��)
T����pԟ!�T\�F��ߔ�P�c�%�&��ͭ�^���˩�F��7��&�����UI��_���
�
36�SG�/�ߍQ���G|,Tml��P�:�=e���χ�؋��y!��[y�z���[?�ܦ�K��he�S�ۦͳ���貲���}
2�����
�������OPz΅�\(7|T됑Q��ӏD>�4���:�Z˸�겯�fj_Ff�-?"T������㺥��7x�*f��e^��0 |أM^\~n2��쎧���-~N4�����8͆?��ۋ$�A��w�����cg�oY�Y�h-�>a�or)�!x�b%r,�Ua��v�iE��fF<=z&����=mY�3���kV�#*��c��=�i��*��]��|n�i�W"Ȃ���� H��\�X��b�"��c;�,"�w<�L�^�o��q��E}Lry,1�./�R Ua���e��k@��y[�x��'$d�0�d��5��Ѐ�fvy�* ��I�� ��(%oT�3�i̚;߉Sl#���WFG��!P��=�x�.xmW7�J����=��/4Y�5�+1s�P��"�fţ;��,����g7R1t�,j�Y�8eq༆��������H�C�œIj�n�.�lBC�dd�Mc��PK���um�^,�{Pf�� �mtp=&$���"�7W4�{����B�k�0�C]�Ǹϒ�XGL�.��ǟS?��#~���F�ׄۡ����R���Wvc L����k䵮��}�%��J/�;�?�Q�n��.����?v�T߁�o�.�Wd�'9�2q��2���7|��OOw[ 93c���[��""�0������f��1�>�H{۲�p�dv7��~/2����l�I�0�-�Q����<y1w1�\Ž�Lb�U�_�c���_�߽�K�l�i�LI�j�Ʒ$�S�X7:��h�V���s���F�0��dI��ۑ��q���5�(����9C����ז{��)�b�9������j�XF���Aø���-�"�F6�et@<(�
�s�t�s�C��3�p��d(Rه0H�ٺ�}v���Dn�32-���n��z�h��訡�L6��_�pfK�9�U_^m;�ݸ�"Y��㖧�#��{b�j3%���ʿ��cM�Cc�S�Y��*�Ie��f{��ȜZ��#������~�YT)�VAMɊ�]B}X��D���o	P1!x(|���'�-�M �U�;�LgP3�
�~�'We����ԍ.�t�Dlv�v��0H��/��[f�q忿�k�6��l~�˯���|*`�����ЊO���J��N   
� ��-W���%�Q��L�h>�~B�((c�0K��*���>~t��s-�]a)-ͽ�6�l��L�q��l�G��¤f~�O��˕g�-��@H����@{���������5��4� /;���|���!�D��!����C�$�)����'B3��>�5�;gX�����PM�M��!���2�.����@I����_��H��b�^X�����z����շ!#��6��~��~p$�N�>�e�ޔ�i� ��+%i�}���1�0�:xܦ���_ՠ�h����z�Aa���(�Ȝ����t=g7\j%�-��x�A�ǶӐ���6�w�����9����%����s�u�7I�iu��,�w��lϵl���>]��[�Q��wB?��1�:W���Sk�%�������d��٥�5���%p	��cg���Rg��B�"0��1�e�L��Cܢ�o�����a�D�(�I�@�)��6.���a̢��r�An7G�Z��S���^ѱ�J K����j�(h���W<��M�
�nyATGl���ʁTJ<���c�IY��+t U�� ���m0����ww�a0�ޚ��9x)U(�Ё��HF�ڔ��@�g`}�3�+no/��Eg�?��y�`B[�'�`�"興�2	x��|�>�"���^M�'��.)Kzw�樞u�����%=�$w?t{5K{��G�!=���L���IJ5�%,4�H�~�m���E�Jل �������yP�o[�`eX��s�N�̫ͷ��9�v��42g/M��G�g��C��+6��p�-�v�t�5d��w�AV"���T�SqG��
;n�3-�'e���e_���".�̞�w;ѯ�] h49�W�`��5�]�(�,sR5�/�F3�#���$���Q��<��k_��?ɡ�(�⼜߉#�v���s[ۗ���־i�R�A`���¢��o�|�v�ė��]d�Fh,�R��Eo c��>�pp�i8twr�q,�ކ����j�������-��;K0�zX��ex���al8���O_�t��ϑIfF?曣x���",m:]� ��6���xu}�`]�Ԑd��r'����T��%$�}(_�Q=��?�0:�<퍎��Ћ�	;=Ip���yP�x�uJ�SE����J��$���g<�a�l����_�(gxř̺���<�N��_���|�z�[�� ����v|�����_� �k�4� �������:ʿg*��'��K/e��L?�ϧ�5>�&�����-���XiЧ}#m�R1�-UY�EO���Z�&w�̡I�@�PI�P!���=��y�����bt�%�:��%�����~m�ֻ���/��g�VUnn�g�4�����MHZ��(��%��	���g��}���ݔa�	D��f�3��_`>�^������IT�M0�i��=��1_�2LW��Q�o*�HA	�I���j\rWU�{G����{�X�(rKښ�Uu��4���,��*�13)Z�HűjF�%�0M/z��v#mX){w�f����7��+��2��
��_�fn�;�;d@B~����?ߨnR�2��k�a�4�y�n�)q(�]p<a��!�'�И{����9�(�8���[��9�₷z>��P�=&2�ouy�v�?��#�(�&Z$%lMo����o��������7M�7��Yn̅V����D#��ϏH�Ĩ�K=�2N�dT���o>D���Ȫ���A��ڦJ|FҰh��\���A�p;���]�6���И�t]��)̴tf���)+Q�;�7�t_L�i]χ����:aFW��o��S5s�>����|�a"���I?yu�~Z�B~�M�{��,G��x�[�ND_kqk�w�%�u-�1�@&�|n�ʅ�e��jl>�Xk�(���PBD�Ed����dl��(���e��ĩY~���(�[V�������^ 썎�:s�����2#������?�iX�8LF݃�����w���X	?ҫF�����/�aQ�DA��Etl�7Ԃ̇���m���b��#��"h�u{ ���73h�?S��ȡ�w�'���Cw��[h�'��3o�0@�N�B"�s���r�����C���޵�dZ`���+�#��}����e�q�8�O��a B׹��>)m�����@��d�:��<���
��|�"��w�u�`�c�s����=�2�ѰV��N:n�&���މw4E�?�fQIn�}_� Z��M؟�X�F	4��B*����0^DU0#�#�v>8��y�um�M��6�Z�W��eT�p1���A�t�� gψnQz�h7�{ơ��ā��f�����s�8�A����:K�Wu�zY�sc�z�Np�$��Y����X�o0�U�=��\�z�>�������ʾ'�q�C�����Sx�ƥ�sk�k|�=n��V[d��R�E��g�횧�]"���d!�[�v�ޝ