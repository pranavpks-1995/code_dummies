3�c'�3��u���Z�wi�.c�F����	��Si҈���`��]������;������q���\'9��Oz�c�����[���T=��vFi(3	�"�Q��J$��2�n��!��2r"��ٷ6!PIy�"���|��kYO�G%�߅D��F��gI�s���-������U������DY_q��>(�ޏ�y ~+�%��~�+5�D%���=Q:�Y�H��/��d�5�<����:H��_|��S�%�ݮ~3��[J�P���Ƈ`�y`�+�a������v�+p<|�n�C��T�R�C"���=�Z��j��'��m�����Ӽ�%K��?�����.(l=�ɩ �1U�������Q���I�C�:%T��%ᔃ[�~f�k�4�e#RV&�8��a:2'S����o��{`�
HB>RLg���h�{X��w�j��o�>�[+Wó��G,!&$^;#X�-#�On9_���i&L���YGUGL�vc�#u#qL��&��8��e�}�ι�wȡޏp���a��f6T����2-SĞ�
PŒ��BG�^䙂 C���f����n�?���xH�4�0�8os]��V����T�w<��8��=l��{��(� d���С|�]!D�fM�H>'�N�z�d�z��}����<��J�p��R"��z�gLad�(<Ȟ%Մ'�8~����r/Z�I��Ss�/Eg���$ڭ�A�b�u���it�ʩ�����v�;�<��KM��r�͓��?+)�eM0�/��k����iʧ+B4��z�7�f����kw�86簱���e���P�����y,�)�O���M�Vx�$�z������P�ao7�]�:���nЋ~J�K�;镩�C�.��y�;�Do}Jٲ�킲���ɝ���v\(��.�����Vä�oP���B�-���6�)X����lۮ���Y�#�l�^��xSR�:-��B�y/g&NF=xJ���P�W�3�r� l����G�I-@�T�a��x!ʻ~ ����P ���m��e��}|�~�$g�wJ���2����1v(�  ��K,]�}�%I�����k*��U�$!�]�@�z�8^�� ����'F��Ou��#�\�����@���F�O�-�psL�v���.��; �p[� @�<���sRx��osB����cbP�g�b�x����ٳl��x�md������i�Ѿ '��w�j�v����\G��'Π��
tY�V�sM�~��ʇQl�ǚ�֤�\;ѧz��O�iݛ��GOF��ZPШ�;�q"��M��,�leRAIB����qi$1���S@�_`U暜U�.�¯W���.ʋ�I�Afe�����yӲS"�ܘ�!��~�ǧ�OS!���d�D�2p.��l�O�ۯ(����,�|M�Yh�gNo��g�j����ӕ�w����B!%�2��b�	�7�R�U�&��FH%����YG��C��������,�ؠ�,	x��D�Я0����>@K��K3_�������Qe\c�����Ty�	2e�)�����u)տ6<���Z|�66��dm�o>_���OPH�mX��`L��R�'\�����xH<����6Ś71a->��?�c��`f�9g`�5\E��%3�M��3�H̠�ſ���x����#n;Ȋi)˨[��p���O�4����vV��逹٪٣:�~z�x�Z[��$F~|���Y'�}p�0{P�.�P�Ǹ�;CHb���U{D�{��'��F2{�_k�8�?9�%�':/Z� 9�\H����)�?�5Ȁ"GY�>���	�!6�%�u�E����~���dT~骪ϊ�}G�L�&h�@�N^/��c�Zb\�>��A�w�KW�:��@dm�֛/��}D�7�;�*���\N�ie~G����\�~�c���y�Y�����.G@u��<��O�`&��l����I���_�C�k����B��	]X��]���6��yK�vW!�}`)� ��</�
��|�y�Q�eߐyf���� �f��tu����'��]�$����b��4~�9�%��s.�*T$£H���n Ґ��
|�H����zSN��+�y�)�) �p�?_���K0a0��v�9D�ݽ��9���3o���嗎�x��X)��_-@ފLy��}	���|�=�h������PtUNr��y�d�Eu�gÉH�#�8�d%�
5�׻'#��<�A?1ۼׁ����n~-ٝ�%�3�EV���%�^Ɣ�G$h��RX����*�/� U�s˓,����.�5����/�`��Џޚ�S6�*�mJ�CC5��E��YH��&�� Z���2��%���:�q��ԅ[��$4@�FH�r�v0՘+�D"�9�� ��8�m�	"7mkk --s�㡩�}���RH4딞�_�r��9k�S#Y�3&CU�M�7A����9�*=<�8�m=�w,�Ԧ��S�7|�����#C>SnW�b��nz*��Ւ>ׄܤ��j��<aB�z�V'�6{�`h�UsG�U���B�;���m�=w�D ���L��n�������!�~4����ũ���E[�*��4�ա�#���
�C�Þ�f?����͞C�^v(��3V���'rK���3� @�4�=��7i�m}�ȹIh'Ԃ0)���a�D�.�BB�	��:���W �xH}i�J�3co�� S�@⋀�z]��h����@����'HV~^I.xq�GOܤ�QsWy��Dʞ�We!^Tؗ���B�Xĕ)Xa����c�s��K�$���� �k�n�A��&����ܑ�*6�r�g�'370izkB#�f=R���sD�&QO�׬q�T�~�`�m��β��.ɔ�S�\~�H��C�W��ؔ={���͹e{H\B�JPi0SD��Y�`���ݾMZȂ��r&�K����a��x��y�S����Z(�ŗEW�᠍�+=9��
�:٦�9>��k+ޯ�z��D-��"�9E_�E8��i���2.a��rlk�D�rմ�p_M!�fֳ���T�s��/u��>�[?��O�or9GO�[_�v��Ԇ����Ǜ���zVf��ɶl�@3���uf�+9s��D�[���}!�б�d�*Æ���Cv*n����T��)�BBv(_�f��R�ɰ��Q>7#���q;Q��5����R��2��M#�`�s��6Z�1�?�ڮi�9�9��1��m`��� to��<fhv����>p|��BK��8U� ("@�W��K��_$P�y(���kK?��#����: ؔ��9׭�#��v�}��"r\(���v��jɽwv��ֱ+���R�أ6��Ŋ"3���{7����}�/����z�`����
�~�^tbg���u$��c!��m����G��y�i_�b��čB�ˈ6���ig�� `�zS�`��+�sS�J�krR+N@��Ls|+�KP���)o�#�U8Frrw�#�0+��V�p�ƝĲVj������8�u���W�JU(��t���J�y+������V��d�B�#bwb����`���ޘ8�h�cv��y�K�����eh�$"��X�_���y���X�z6��-֏uدr�T9�Qܙ/rh�k�4 �[����("E�4��m�������5�`�����0���f����+!��-<��n�/O�cc�Xk~����).��U+ ����Bu���#U�Ͷ/��E�h��\)��dԬ�[}v#�/]��ڦ�V�0���&�bϦ5Y����L�!��r �x�u�,Y�r�� S+��yN�
�i�!l^�d{� �dؽ��K}���8��O�j|����d���K�ed�,\G�b��t�$�Y�H����6��R�O:��%���T+.xoݭꔥ��?���o|�:u���U&Nߘ�E�`��5m�iy�`S��*��3JU5%J:-�X�B���W�$I���i��jlq�h�ئ��ko��!&�cǛJT͕(ڛ� �[\��&�B���?ٳ�0/�0a���3�%�F~ �O���j1)<3��d�3��mޒkn��Cݪ-��|N�o(��z-{�����9��#*�p�����ث���	��p]�wZ�A���C�O:�+��H�{�-����*���=���J��3>�j�����kX �(����<����~ڬ�[!��F(P�+�JAj���1�u���|�����_Fw:�wq�U���;�(�������q����j }�2E�d� F��D}Z���ݜ�uB��g�v�ܾ�|��G���4bN�Ƀ[���*|�+���2��:��v�6�wF��Ov;��:��P��]�mO{�fAkI��o�)X�)����<Q�d�an� sO	�v5�u��[+�l�7IƏ�j*�O5�ȵO9TC�Di�֭��������"g�;��=�ݚ��_�%S�5s�<|#�L��i:R�"�
ڼ�1���Ƈ\us�̞�t�]}[�v�( Cy�G@U�|����L[T�w���FPzF��%% o�Fd��"�*�g��ci̕R_z�9�h����1�}a����Za������n����Y���?"}�Gj�ټҙt�j�
Y�(�	0M7x��y�lW�3;BQ�%�~���M&+Lj���F���� ��j���z�KN�7Ӧ¡20����<���.$��?Hq�����q��U��n۪�N�u�����[",�.Nk���ZcYlI��|gЯg��A����Җ��� �'��uG�i���ѳ�L�'e=�4����d���(;>�H%����}�Q=9�"難t=RK�):�D�h�*�tF�T��i�f��-��8I����k�	�}
��In`�����Z5߲~��Mlk��?�Th�X���C�D�=�Ţ��b~\ۂuM�Isg{�?�	��(�DH�1awY��Qh��������"x|��(~��s,F�(07b�L�R��j|�]`*�/�WM�u�d,���:!�������9��Yo��s`��3�a,ay��a������.�B#�
h��r��/r��W^w�~l��7�rU��c��wgE��ͼ��=��<HoU�x��]�uƅ���7Y!���֒2�pN���V