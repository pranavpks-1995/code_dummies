`(t(/ =(��[��Rv>\�$��������6���XD<��r�-�"?3����I.��h�p��p�qR��x��iQ�Gy����۲����ɤ��������x��~�t,ų���C�/ �`�lيN�h�����~듰����ֵ�'�,͂jyf�d] ƶ}�^�+����կ12��LR���W�f��e�A��=4?h���b��Âd)����fG���@̅�*�E��+��dE��`Q�}�7�d�"ai��,L�vko�Ks�C�:��Z5P�yzH�{��*H`���X�f&�����v����R�_zvt暘Ώ9vdN�@e\Lq{
��P,���Cݳ�Ƞ�;p5A2\ 4�vn6�ࠜ�F�`P]��?,'�Q͐o��R�x�Tӷ8���\�1FoR�e�Yj��+�V+@�{��We���j�d�w���i����]Q�-蝥��()˭�s�%�RN��� ���'��I#qԟ~����'��A�|f�O+y���1��ѹ��0y<W���1G_�&���n���{�:�����ב�+�S:0��9:���e���Gi	̒>�M�B�PΦ,PB�D���x����/y�L�7��8�X}�KM�z.�|��*�#�o���L�$�*��dY��������Y������c���TͰ�s�`445�F)o?=|+���-#cMe1N���&r�.'n�	��w�$��ϯ^�@6�v�[�כ�����'i�$?�h8m�  B,Z���WWS��<������͢��s'�/�a�h�a{]��K`����1�kF��3B�?a���zjb��h-8>$k����%t����uř����~ۋ�X����Lf��p��=,ϼP�d�����g�Ee���Dwd�+�yJS�g(V�l�R, �,��%E�RӬ�k�v���Z�����Iwu��#��AA5u��(7��W��12���������S��&�2�I514�ϭ-����R${r�i�xM�3��y5��\ø'M��
ˤ��:�����l�![�\����h
�Vq$1Q��||�g��a떂c�2Fs�E5}�Ǆ�|
�LFdZ�*R¨'��;`YS�ЫC��L�}c~�{_�o� �i�"��v�fen9�Ê^ ӓ�����Df為����é��]ʝNkoL���5{�SUv|�i���]���Z��$�q�<+������ʂv�KS��N�% ����q��B��<!,mTS��������uP.5JcM�E�a�,8��l8���!�߶t�͉��<[�[��/�X�(qoG�$�J9bz��=(]x��NId9�툻�!qL|�7g��R�5;Z�SOJLK:��Y8c��]����sID�^l�`��������Q�g�9Q3�l���îL"9�hU����wJ��� �ߨ\��{�|��}T��*�k֘���1��������C�A-�9�
p��OP��Ӎ�x/�_PF�+Hy
C�r���#{F~��Cbu0�j�(��{��d_;m�w�l}�ɫ �E���Q&dÈ�s�:G��K(�V�Anu���n���}�l�2y��~_�E��3�-�et�Ń:ge�m2>X��I�6��F�j�5���7
�R��>����-B�4��6��?��סys(��G�X/g���̷�}$�T�zף�)���C����i1�i~�����蟭�����+�R'�ak<��a�_��{'�����|��ON����qLXH�K;�z`���0���v�yHJ
8nPIZ[��,��%��+;;%�q��9�
0�ƂM�Y>�F��gHف��;�=Ӗ��<#����k��$�=��k��nkEôm^�%¨��(�ϖŴ�&��h�D�-a�&�_�T:��h잯\�U��.���ĩ����ԤSI 콚,%_ ��?��|a����S�6N�b�8u��u0�GvS�GgIr:�����;yk�/w���vh��vl?�8�E�$Y�+a	iZ��+��	H�iy� E.],Y��o�&�F��[��X��渷�����5:E���5	��W�>���N�˪.��&��W���mZ��D[V��,�� gXƷ�{T�nH�6�M"��Y��!��ر��}�2�&�~�L;��ґu��z�ys)�d�y��C�F�S}T� @�w[y=͏Q�DV�k��4ع�����K�I��mj��qwr��Y��U�YI��l��o�vd��@��ү���Ţs������$�{&���:r�ǲ��l&�=�;LW�06P�(b�Q���3�VD���#����Ā��P�#M�a��I䦌�6j�oY�?�L67�XvN�@:�P�Ap�0�B��n���D��~����~k��O�
�O1N�\M�KN�<�5��
�3�	��&���6��I����y�M���5�Q6��!�+�=��� �M��l�ط��27F�D�����O�YJ��Ǖ<�� �ʂ1o�X��Z��k������Y�jʣ;^v�Bh���9Gt�V$�����*0~Já�
�3��C��n:d��4����q��CQ�\�&�2|񞡋��ϾLKg[��\6�D���h��'��	��0�Q�㎺��;�'2���F���=���ۣ+x!��.�[\%��q�ؘ/ʫ$G=o�ǾN�#\��v�k����l�uJ$�I4MR��#��o�a
���
Á� �J}ĥRP�e���[89&Z� v�σ�(D���Z�t&�i�;����k1+J�D�`$~��\�S�0�{�d�MQ��b���5r�3Ш�#;�:���'�Q��|�um���ug�6:���N�kᵹ����w��\�A�B���b���2����9+�� ���4V��'�Bu�N�_����oB�6�{�dQ�n`=�W�T���}��o���4[��mo��pus��hΓ0�۸�'I���sAH�ꕼ�1�VW�vwd��#�-��*m.8��E�4(C1�[tC�����Kr��i0d���=��2�A���O��]�H��ڊ���������+����<�����=�p�R�G����n���,K}�fW��@���QX�i}>�C�M�sW�#=�T����̲��l�젧��%�XY`��	*H�0���v�d0��xCVr�B�"�� ����^�zg,/G�z�����=X��۞��] ��Ob��*�E�g:�	�[�iZ�2�R�J���M�(�w<�Jnf�uH��+�a�G��7�3����I�>R����!���M_0���6`��M�_~j�h�h���3EȘ �0y"������<UN������n�T�ܑ4�V&Ƹ�$���;�$d
��#�ɇKi`��x1�07���M�oI� 9B�I�𘩛��m�~-F��J�G/�}Mz���
>��4F/��A��Kh��N�S#3��l~�;�$�-�c�i��'��\$iSY	g�*0�lQ;Á3c{�[n��i��pL�YR���}/���l�;�<q��do�}.�p2�<�^}�l��;���9�D���8cg6��W���9ϗKe�j9�v�5с�j	�����"r�uJ[�Psv���n#*�z�_�����v��C���m'? IL�����	=Ίg/<�)x��e���F�t�J�`>�Ā,�u�r5�x��:-NĐ������n�5K��Z��x��G<�-���J �h��\�Ӽh��?@�T�� d4�}�5v��c���l���w�#��N�����p�W��e؝��]��4L���{����P��h�emM��]|'=��j�R�
j�Ew���F��HІ��O�K�R)��vˌ��s�k��f�F��sMc�\���c1���ώE��� �gu�N˨���Ho��s����(}��x�ލ�d2*�x�~.��K���@�0�Uo��~<���������l�t*V��6�tc�(3�L� n�O��ׯ���Q�
�>��"Չ�"�zdy2ۯ��Ai7O��)�O̧#�����K�Yg-ש	�/c�2���o��K�&:��C&3+��c��M�l�́���DY�
[,~��3�%���R9~��Х�d�Gv>(��d@�d�ӮV:�WQ>C=E%eP��dD=zT^+�~pg��4��$64�}�W���>�[�����r���ϬV�踹&���_'W�s��q�n` ۫�t.���~;��'4&05i�V'r�ǈ�Lpa<�h�Gm�v� �=fy�N`�QW�*%����Qn��� ���
��op�+t�mx��J��.G�c��[� �,�*r�Q��-\P-;���;���0�GzHc����<�

�N��5�D��;�E{M��K�Jڧ�� �+���;G��q��iÕ�-tz���u���R�~2`�/0.\:�g�c�d݌���l	B��u���nW�X6ثGx��+@`�͘)e8�d��H�Pm��8�a�������</�O���.�����vw��
� �q���?:W��ZG[&"��I�=  	�'R��c��s:1ĂaHB�8�/c'{M�:�ffV<u7+���d����<C�ziE�ǫ��n^Qj�5W��\
ޥX'GWV.=�%@���1�Q�9Q�˯�Ѹ�X��B.|�]�������DǍp"֊��C��s1���'z��lt��Rj�cof?���2�E�����0�Z�u�+ۻ��hLS��T�d���z����X�>����Y�S�q��k0�H�S��Bk�#0�lV�o�t�j;�#3��ڧ���)�{ϥ<��j�r5w��j�$���t9�@���(��?6�{N�c�:q��׋�/�[>|O#��Em`�W���1@iKT�s\1Y��^�B���`ZX�=��o�t�0��{�N�i�#�Ot/D�V[`���c����~ ���J���.��y�Vf��|ω���19�N,�@)��dz4,���l�kȈ�f��4���Imx�1�M�!�5��lb�4cK� q�����ܖ�-�#�����v��+Z�r&烠���l��G�G�Q��\G� N���~�������zq�"<0����K-yhiŅ�����Џ�&>u(^�WV�yV��ߔ�<�i��d�)�В����$��tp�ia h��#DF�z���?|/�rE�X���^r��A��~���c������G��$�Z�$Qϯպ/n�}�W����w7s�g��'Xe���=srX<
�Ns^���GP"����>V�UAԙ.�JO�sj�sC� N"� F��m�a�e�d>��#��C�� �|��g�:��w���-�~�Y���vU�N*�N�}l���S��.q�[E���;n����9
�n2yx�/uz*{���iK��)Jg@�b��%ss8xoCU�w���Uuv][�-��ؓ)0�M	F���"�92��콺jh�%�Ǖ^�V�fزr�9lC��ǛA���\n|O���b��bW'�N1y��H& �A��l�"�Vˢ�5��p4i�x�\�[�b�m�
�������d�0�
��HڔB�e�@������y�^J<&�K�*���-Ϗ��br���qқ��=�[��e�Mބ�;��X�x�p�l��/1�h�v�V��~���XՉn����?���?*n���q��6�Kݲ�\��w��6[)ige=i����C���a��� !��ğ���Y���:�*�d_x#�C�^��.�-���hzvj�?��`ͅ��>��������٬��dur^�7d�P�R�r0�w��PWHW)7���o ��LK݁�CK��8�g��������K��&���_���*e/�UP��	��c��Z�	�2�qՐ/��R:�ޡ�������P�_��93����a�9�u�����U^��
2!k��}R��-��'�J��P��*x�x��*�gV�$�u�l����Y*u��_��F��h~rT�� �w�$���_a[���~��u�XL��fb�`8��_�s;�*@�d��P��x7�p�k!-�@�h��
����lm'�B]��?���z�������W����M��ɤ͛��!`f��Ƥ���1��3��r}�e���<2�Q)H��9Q�{}�͕ 6�?h=�u��1�w.7T��V�����'�XW~��D�%����L,�%�%�^b�����bh������Ҷ4��)�+���,:�Ā��no�P�~������ཟ\�LGH�-?6�
��R��u��t8o�S������/}����I�=y���}�����g��n e��{���֏@��,�s�p�K:;5w�����]�>u��D﫬�9�O{�i�P��I��x.�[l�0� ����W�;P�\徺+|���E<.C�¨�l:�Z��B;�7��ft����r�~-@���H=y	俧�X��6�G�iD�J0u��ܧ5�F���;`,������XQ����ԯU�4W�^���w���4�U�mN)���[��SR��s��J�>�A�@k}�#ѿ��a0���A�<����ҕ7��r�gr��&�6���C����Ͻ�	q�0k���3;-Td&�A��I�3r9����1b~��q�3T��܀T��� �@�s�����T�g�ۭT*�<�*��Ek��$��֜2g�`��6���Ć��9;�`�(j���|�[�X^��)�Z<�\z�AXW`A�5��`,^�%긐Y"�j~�XP�!����K6dQ��&{=h� �	�<uwc�����X��@N��K,�����^k����@��d)�E����!�s��2�[��@�Eہ�  � �F�U�&��c��:��6L���7���C�
����w��]>8���Z|a�͏��Gm Y��y��B�3�J��,���DRW�IO>�i��&4㞁�������٦Q��Y)��x�Dhb$���Y/�v�+���q�%e�M�EL|�_�>x�_lH��h����_$k�x����f�Eq�N�f��}�'�R�϶�4��C�������t�O�`���S`-p�[%NR+�F���)kr����b�@��n�XV���Y�<�[���X�EDb���I�!���H�Y!.�ZS������7ZutIO�CHB����W�W�ʃ��'r����F�/��j �_�2E �Adf@G6����K�F�+M&J&��bV+�	���I ,��-3BF��I�j��@ ����Wc�{��>Ě�������NEm�a�]���d�,�:���U��2İǼ2hQ�����D��>���Xe~Ѓd��p�~��j�M�(���H��h��v� ����-F��:]?"b�ti�^e>d�Y�Z��<D��2+)�������R�j.!5m#K޷�(fW�9@�w2��t��� ����	-�`��St{@�C�I�����w��U=kꚳ�H�Ƚ{w7���v�m(/�v�����@{� e{C�ڪ���I��w�J���k�Q�	O p�=1\�Cz����Z+���٤��i���(��C��<�Bu�~�s��Z#{�9(�f�kD��2{G�w�9ᛧ�V0S�r������h���J�����0_q}މRu�b���L<v�yɈ ��a�����C��ԉ�NB�ͳ14����ʌr��=�&��[�xDz6����r!�v�͊0�辕B3q���n�6|�qCj�'#�nMT(�oz�Ɔ�2�신��{R������祬�i77�'����BQ�4����Z7�2z�!����3����S~�K���{��T�B�	_���`>H멻 �>Jz���o!^��=��Is��ZS��v	n/9U_�b�������X�ţf�D_�(6y�u��S�Qd���M�esǜ~���z4��v�S8h�q�t0�����y�G����c��o����T�\!�#��Xz}�7�.�{4��f�ZN��\��[٬��o�G�(��-�����r��ر7jI�sƖ��6�`=ku�Ǚ������$��;���>�ibwj����E/D�l\�ˌI�2�V� ͻ�-