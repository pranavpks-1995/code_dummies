V�f�iK(��OU���S��J�����)YEF(U� dmM6�mp��w2㸭�!���|���T��#�0R�9�H���So�0v�*��0+3�y͙��w����J�T&��_���T5=H��0���|tyK�o�!���$뇀x�=K��c�28�Pcڔ@_����c��|�)dg_i�	X��o9�y�Z���W����.��۟�212c�`�:M���M����~9�U&���Q�#��6O��m�kq����h��u�̹�����6��j)h� �E��V���,�Fɧi,�� ͝�:��Y:۳!Ψ����c,�E�;��{��HL��'i��xl;�?׹ȭ��yX/���u�~l�)��"�{�7۽w�����au��]���Pu�]�!y���c���Vd�\�Fh7�A�|����C������~lÚ�
�Ծ�� [�6��������T�U9�a�K2���q�"ԇ�m��N�~�n�&��] �u{g��y�d��,ז>�g�2�o�����"��cR!�e��<q��1,�ƸKA�[�>�f�%��%�б�/XTᩀ�(�hЄ��&�܏3�^�WnCǴhx:%hvp��K��֊�k���.���3��l=�w'E �e-]7��drs���k�j
TB�7o-�|���E3]M�����`b"j1�qk9GX�QKk�J�d�V@j4a�pi�5@��߇z�\<�fh�Q��P��L��9����B)�   ! ��-�����L����RZļ
^�19l��LX/�P[9=�0k�3�������¬.�����~��HKssYe��[�/d��q<�q�^, �����CGbAFA;��cDy���E��+{�9��W�"��� pd�H�>�kX��&M��C?�����]l��q�`
�������} ??7�E��QD����(��e�̓��e#UjP$bG����>���YӒ�� ��Ώ�9��!�`Ǧ8�2�w�j�,$qټ!1J��yJAD�k�������h5���Aў�Y�MQ��SYL�m�=એ6�	~w�YTuO7b=�"�	f�B���&� �i2i���x~4�'!�Ј��3��\�Z���W5%���نd\/U����Ƹp���־>%M�^W3�^�s~�N�n(�WA�4�B7����}�~�ͪ����;6� j�PF�`��-5�L����6��"�Y�j��G&D���zA1S��x��VV��f��DWV�xɖ>�����������424�%��c������9�%H���i��t��Q��   Р�U��C���J��e��a�C�J��h��9��.NK�]�XkZ��[IF�!����n(��#�G0��� ��v�v��2�����d0����S��w�P<WMH�cs���Bd7C�s�)�)-k��B�������dg3n7Kw�w�˳Z�n�00{*k���4�,��qy��S(��Ӄ�F����q�<F��9%3�Z�s:��v�R ʩy�
Ʌ��1�#��a/V�<��f{A%�a��[-C�����|ijf 0�C�A:Ʈ���.�-x���ʊ/t�,�&������=۩�da���
Y�n�P�!��Oq���������f���yy�`-�,{���`������<��������>;pp�����  ͈l�e����쾆�����2�8��7���g��|O�7�� Q.T!��sf�6�.������G8,()�~�~��mx��U/5�ŦK��;�u�~�ˑ�JC�H���N�[.DHcqzӰ���h�����P*[%:)��[pEr=h�\��`{e�u����l �-��X%��1�F̗��)�Q�j�����~���R �C�}���M����0�Y��.�e�9�v2�
�C~b����k��a��%�(����X����y�rE/������������mw����9�l�����Փ�?��A�3Y;��fX�:���ַXq�mh�GI�.1Wi���ۗo`Wg ��9�=:�ݸ��\�]�ft���>�Y�{d4ԕr�[*�	<~����]c�074%�z��v�%���h�IG���M��[gg=y)ٹ�G�2���у�l>Y����KӂN������ ��b��jd^�K��!�Ъb`�F� �.��:Ļ�kI�Cpӳ�i�{c=ʦ�c�,��F�ص�iB*�VB�Z�D�r�B�[|�]L����A�޵qŞ�4T�K��*��k�3^k5NϻJ�d��!���0�?'��Q$��5�;eSsC��M�^S.u=���}�)�S�OjEy�+�G������N�f���殅9���EF�XMIe�tR5b�)5/G����䍇�FJDG���E�&W}+�Z�:t�Krt'q��P�!�?��`��lK�釜A��6e���d�E�)�54-�i���W�uo-o�:/+��@�>�\�>&h*�=�+R��;4n�BX|��llb?=���ª�~4��>����E\��X���òH�n?󻅖�J߅7�c��K��^��Ҩ\���UA���A�����d~1M���nۭ����j?���
�� "g3xjC�b�g�ԋ}{�"�8����*�P�xQ�g?Kύb>aL��x��- |@�*�

����}�mۙVg��:O�������t��5����͍�  �d��`S��Jgiؑ$����g{��Y�̤�T�$�H~���B��o3u�Og�`�X։�J����^���\T���f�lu�f��n,T������J����&�����п���ʔ���4��Ѩ!|�^�f$A���{c*(�����h�W=�gea5���F	~e���}*(xb���'3�V?�0��WJ-����� ;��@E;���H��e�=N��vh��~փH�\�%�+ Q���t ����hG�*dp��#PP^���bo5
�.W�Fa@ey�6�>%�!����w���'���[��)o2ӕ����b&��7qFx�\�`��j���zcB�w/��S73>4��}���0��!�_�� \��$�8�{1P��Üϋ�i���&�W!��Z��4kx�����%��*��&�`�������A���̲�L!�p�͡��^	�K�=�]qF`;��[cL1��
��\�>{sbO�/�E��:W�AԤ�ޖZ	�4��I���CxB`���#�-��A��@���T�V��e�t��~R�~؏$�k�o�9�UW�'+XP�s�|��`0%��9�����~����]I54�&�e�5��\tЋ�c㩑�@�/�Y1�Rf�����D��lm�?fI�.���|�M�1�S��i�L��#�~��l����厃-�GyT'��;�V���OcZ��G?��_nԕ	�"F�^fE೓�؆&�^~1�36*�ȓi'ϧ��P*���~e����Ů��9ּ5���@ C����zـ��)�}���g:0������/%=U!�D��`�E�Y������A�m�qRM��ۆ���KwH8O��G���h<R�ˊn����-��<�Rb�����{�c��,Y�����߭t%~��dy��`�?�0�"����Ax$�y���c��6�):�65#�%OC)Pu%QK����j&�U����Z6�@��涕�"�oISy����c���6v��6�șI;���V���k.	-]�8?;�q��.�H�e񨝢@�?AO���+�7f,���e*읐�s.��Qk��3�n�(���ˤ�4=* ��~�v�O���Ps��5�'#x{��Υ�'v�9���E+L����k�i���9�[8�C�����$��pg�ҫ�����hp�zr�uw[��/�\ы����R|�}�A}-<BV�q���[}/��W���>�� ������ũ(���gY}�>4�v4��o�l ��)��FD�%ڧ�L��ڥ߰�Y]�`�;m3��)����o�y;����Z%�K�(�jS'��Z�1��c�ݓJ�U/���WZ�}�]Y:?13)�#�<����g;�pja/���I��S�J�1�bp�HqT�p�LC ���.)�
���<n�'�A�\Ԣ9����Ly]Q��������b/��vnʉ@�`2��穙�毪<���l�p��G�'��Ĉ!<�u=��S,ԨF���[�J�z�w�T㲚���WX9_c�2O��Fj����V6����w�~�b��������~���j�M�+���?��:������Q�}�u���FC��l���3���%2�B3�;�@�Fp c���+����6���\�*/�+�\�R��W����>F+�$F��D'��K��w����S�)J�o��[���4��)����A�?i�~*GB��Z��酵�a��ǵO��ZՉ7]���6��lg'�¢iO�����80cg0��������4H�!�Փ��s�a�%XRmU�x�
�4˱�����@IUN�Fv8�Ns��n�X~�FW��5��ݧ#Mb�:�ôՔ���(�F4M��@ߥs�����v��` E����NT��mj�Q-u�@�p�n�%̪9K�˿]��s�׉O��S�$��i@8~�{���ӯ^O��%�
�NC�ZSx��2������B��֞F���Udn�¸�6Tv}�����z��n����T����/�Xj�p���@M��ϻ��Os�_X����iɪ��oX�ڸ{v���T+k7
��D~�x8vx��8�����M����"`�[���e�Sd�c߰�s�>4�pCB���Z��[�z3���	�;��[��^������;��9���&��xj$��:�8�>��=�щ�J��LL�FA�uUyr�Ց!yT�K����3]�ZF���s=��<@+�3�T���7��C�4>{�v0�G�Q��p�^p�nUؖ�`�(]���5����C�S�}�+8�Sώ(V��j�#��V�]V$��ʣ%��c���_�l_�ӛC�ӆ�L�0���ၐFh����ç1��¾`)��.��N�)���A+%[!��r�
{-r2�-�"���}S��c2Y�b{&���n���[B�l�~����-hG�a��X�)��lR\G#Z�̬���Bk<$F����}����g.��Y�w yc���W?m���R���3!p��|S��_�M�?5�{�+��hq�A�[���V��3�Z�(-�U��7?�O�;��\�%�
eǟ�}���LA3�\�=hN	.�`���k7MA3���ɶ_��vm���[k�(~���!K��g�f�i�
���̟ۜ��t!q�Aj��}1��X��������l�m�������lfЛ�\��ŤN�wհ�7�>�Aqw�3F�(�Э]�m�Q�=�c?u�X�4y�h�X=WPV�`�5^/���3�u���NIb�;���>�Q����;�eS�*�a_����/���k�3�Ȋ�>��pY��Sr��0;�.��`�:�sT�vn/y�W<�j��������i����Dǁ�  ��B%R��c�����|K#��������#%^΍��畂�k'����T�U�#��Y��q`�PR�~EG'���"щ%,�V��S�[(��(S��"ޓTH���v?����S쬠N#Vw��v�|�[Og'�����4wT�)��I�Dp�����P�
����Sl\z�@�1�*��ҭ?X@Vi�ʄ��U��:��8U�{�ƾX;p���Q0��`����.a�y�=�MS���a^-(��"xĦ�C�]H@�6
\0^Ԭ!�#V��{���И��D�Ϭ|�Сk+�q]��Ҡ���+�+V�4Q2�}v�{�M���E�5t�ԡ�������q'�4���ޢ�j#Ƙ��0����|ަ�#7W.le�H-�Q$������IG�Z	�P7��@&��1�K����H�A�ЯvF���.>̩�_\eו{���H�Ԯ)����s��@G��[%a ��J�rJe�����iZ��t{ �0r	,�nå�&��㹢��7jRԮ������L��u�8ҡ"��C̬�ۏ5�F�ߋ�%��M",���g�Z����k;����Lǿ��d
Cx6E�R|���MUP��X1�i���н�a��QJ�C�y�r���C��t841��(�3�5)4��\ �k%���|]l�CT��wǃ�b��}·) e i�*�B�AIV��DH��
����Sb痿c���w��:ș�~y���?1��'�����\�Т�N�r�@ПU�+}=V�h��̌ �ߌ��2�,��"$KR��b4RR�[�L����J�k�� zBӅ��t^>�M0�	��N��9u�>Wz�43�%�0Ï�r���4aO�=ֽ?�uǀ\�X�:�Gz�����ruSl�[B�/؄��+����O�����c��W�[�Z���b�*8:Y6b!ˎ�����RKMG�dewM�5s�|�����Own��s�`!�h
�m%Vv��z^a�5A�V�OљE25�H�T�.i:�^(b�2�Y4�$��i�1t��Ns���;��|�2������*�\7�)�Ld�����y< ?���A�I��3��z������B\�,Sx�Q��s�������na�u;��)�*�T��'�z�#����ad�� ���3��7TK􃂻�L��eS�XH��!�O4㯍�a��l:��.��{fڠ��X��r8�:8�N�<�c�ΣB�b   �&���,t`���ӈ� �r����_�`��M�[��¾>��*ʱЄg�F��̃��&��3�^�/��T�3�e�A�� �d�q��LX��\b�&c0o��L�6q�8��1 �t�^!]N5U��#dM�*ˍs��^��6�1ϯp�e�2r�	��.�
���nqC�%������ɨt� i�q�ъ�\�$ff��M�@mH�/IcN9ȏ������A|8X��_DB۶PT_�+`�r��*���1��H�,gt���{T�|l���K�pzqjeji�E}}@J;׶�V�姗��Ȯ��`��N �����4��e�o.,5��^��N����P�o�_�FP>�� ĉ����C�������f�5V��Q��xB�Wy8&�+rm�F����G|^@���z������~����/@G�����G�>G�����u���jnX{+ Y ;2Y��P9���@�}H|O�a����6��`�
��ࠪN ��63]SV��4E<��O�P���u��Nr�@�y�A���   � �b-W����R����XJ����Gu���8@�2#dUw^����=���K=��h��)c�'��?"�/j#AXS�>�G�@��߮v����ʙY��Y�>�MEr�!>|��&���6�x�DUׄ3Q��|�� rD�;��7���FH�I��h}\�8� �94��E;��&us��᾵h["�Mz�Tmt�,72��`7 �ѹ=��'cN�����i��gd��݃�f�������8��H,�����!���Z�+?�\��Asn���O��al���i��[��m V���(@MPu��%�<n:��4/R�ȳL}zs;���Uv@�o�S_7Q�̴M��1�/GH%h�j��%�\��?H��t���R5��b���P28���tiǺ�]��8 �����m��b�ZL��n��Eb�_��������!���b�)�4� @�U���D!
�/��87gH�'cx�b�q%�ʌA��Z�J��u|>��d�\o7T� P���:[�;��@�����ғ�nݚ�e��ŀ�/MSQ�B-z��t�"�����4�h�o��QO�!  �D!p�� \���<���oՔ��Ӻ��    �!����/B@� \�5��/�v�o+ڻ˲��X%1?⍷N,�(�S�@8�����(�0����%zS�"��Ġ�w�)S�p`�v~43�j|���C�BN�9&�m�)P�;��U�#���Cz ��n�cI�V�]#7T�'�;~��U�    !����& ���"� @�)��H�7��qy���;���}uRѻ1�	<s	������Z�@����4v>�خ�����0�X6�� �� �v�񽰭�ug۪������+�������u�s]D
A� ��S��>���`Y\��UqP���<�?4�v�j�1�M�B
��ճ@`L`!��ĥ6��h1  ��T�/ [r�󖴜>�ɰ�w��uo�w����Ց����ۗ��ll9����}�w��4��LI1L}#���-���ui#&�R����&-3<���l�
r���x� �߾�� M���]-��rmF�]#T�U(q�v|�@    !���#���D�	��-Gb\k�B�X�`sd�Z��Z4�O/w#�L۝	�;�'ǧ.`{�� "��`t��̒) >�Ķ.�R{���Yo!.S�FF�5C��I�4�(�����>p�IS(]� (�&D�� t�7��j}=o��\@`  p!���`��h!*� 7`i`'�*�a��U��Z�YDp>7���L	� ��qHI�}���#1��������tB��QȈ\Yˢ�I n��\���͹��?���KKLϞ"?�)δwFѩ�	@��8 
��ӷ�����˵��9V�m� `   ` p!����a!  *-M����|W=]jz̙�̱,Ås�p	�jؘ��E�!*rO ���bL���Y5* g�5�5�P
�&fqj�x߱��|k,-=_W5-��CC�:al�P�^�;��!<���O�4+#���͖?x �!�!{
��]�{� B�O����ϑ� 0!����$��HAV +��`��!��DD�+<��l�~B�����j���S�p�U�U��$�M8<!0b�1B��	_8��´>]�w'?��X;-����� 4a܄D��x�S�MDu��uE5���M0]Ϫ�~�L@%Ta <��uz�Hp[^�����n�   �K���   ����UW�C���v@r[*#�:�s�`�'iL��}�6�<rش;�}�'�$R�N��6��,�XʚWޱ��͚q��z��<����o���+�W��63V-�m'�"�ˍ�2���y|�;K V:9�Y⛤��[�����N𯒄�I0�RdG���E7��SgD|����$�Lf�C�^ns��r�+���t�|�喝�1Y�p lW��p%O9]d�і�0�����W���1GXP7�p�&O�;��5P�����͍���y鑇���,B �`]�vC՞ ��F�����4����Tx��K��]������̻O��1�E���긚�g��V½���S�o�Fo`\M��"]*1:� �:L��u��s�uw��~g}�	���j��S