KyEYݒ+�~���B#�҃�vj��5,`��c�ø�?��5`�:Y�q�8K�5�a����ھ���h��)n�w���9���g���`��O�C��L�GAp�-~��T.��3�Vc%�Z��ҥ �R�$�V��E߀[XZ.h'���]�q���r�@]��v�2/)�U~����O��.`����58�3ې��X����uN;�D���$>����j�=To#C�nE�t���S��k��F���q�r�#:6��+�y!��Ad�3	�]�u��^��s6�78���̮@�iVpڌ�69�N�S�c�~kqDw��-������������<�=��F�����m�����W)��Mg��{iࢯwzk�9�b��U�^^���k|��n���]����:�6n�1��'���|<3�B�G�������qI�"��6t~9��ж�hd�w�vH�k��>sf��q�ʏ�QfF ��� Y�7��!K�f�,�����cA�r��ߥQYY�9��ňT�L"��R���cH;�Ψ�*h����;�;��)�-fI݀c��y{�N�� -C�/o���?�7m�?�Z���]/|��-�o�<�n8ڨ^8+��7��P�Xԋ'X}0��{����9��-����Π�o���A�rUL�@�+��tz9�\G|�'��7=���-�:�%�2�zp�e�\� pG��w�~x��p{��QO�4��3����"�LI:���]ɃY1���	n��늾����n,�E�(��EI�h���f��u�t��jD0 �[4�+OW��������╄��MN� ��J�Ƒ��*B���*sM�/�{�)�ᗰ���#	̿�b�����m��,6RV�2K�k��K��f6��tش��wA M= C��~�,�N�I�x�\μ����mb1a�oRDz�Q&���Q��5'�8�|�I�Yo�+D~�\=Ych�A�cC�h�,��A���g�*�bb�|��m ��̦�J�j4��!G;y�K�7Iu�x��;{��o.�b��GV�km_�2�����R�J�냩%`��G�Pl�6l%�����4p[�����vG+(ۮ �Y�vwbfX_�nH����>_[��
�4������B�V�?�s��yԞZ^�`m��}��P��o��T��'���"���������Ay33��m^c�8>Bz2
��;���)k+�\G�Q��G �-i���]+�(ʍ�h43PO�h��h۞�� n�L��1��0��
O#r��΄�'� ��5{j�+��~~F$�Ĳ|���s�I�>�i�+Ɉ|A��ppl93b��U���{%����z[:����w�t��:h)��Ai׺�ĵ^��@�-�|Ѩv,��[�~�<�HQ$�j��Q��؈�aX�g��n8�;����>\�z��y�3��!�Â`���V�dV�J0�7'��@Y���+��R��bF�Wz�#���vwvsW�a��;� ��;�a�TK��$����������>(G!���u|] @Y���~���1���i��ɬ$�$0�7��5 Dz�5��3s3�p��7� y_�n��)�l��:8oaa��V(Y.�s��'1�Cb��P�4�&^�
ee�/��{7��%�'��N�v?�jifX%<�(A��n�L�H�L���VqPm����`B��MF�7p�KlUf �ڣ������6$�E3Z�2��ц	��ɂ�FI�y#���f�l��ea�V�����:�|�J�D�'����OL�p82������J���.�['n6yw�ֈU!�����cB���|�J�`o5�l��
�ou�-.���R�l*#5r=V�!��9_�;�{q��KL�T�7~�-�+���o#�@$m��7s��C5#~#.��.��/��M����t�lLh����c�#��a����C��L��5�/�r��z=�x�e�p݉ם�"��
��l�|���*�-_�d�d��p�Ov�Isk	i�!m����꡸s��)q!Om:�?|��ϼ��0��d7�����k8��G�#�qY�5c�͒k�"7�4�ҭ�op6��������гt�G�|XS��1��,2d�[;��N��!�p>����Yd��tD�䣪1E�_u�:a%���a ���V����f����j&.�V��H��j���{SF*9q�X�d	�'$W�7bp��x�!�	�D�M��o� P�5��M�j���?�c�i� ����Q�8� �J�`��چ�2��!��bQRJ�'Li$�����O�3��� �<0��?}�� �JoJ(S�T�dq5�@��9�x�Jn�J�bŴ�-B���*aԞ���� �� �J��:L����}W�t����P�!�mA3S�8��\�qШ�ԹL�{<����Q�yqI��<��?dRr=C���L����'M,* إ�./����_Vm }�Qٜ��S���)a�u�>&���8f�pe_9�ޚ� 1�AH6�K<g&��ӗ�������y�ȗ3<ջ�
cD���u�Z���p� =�9��������kP�+2�Q>�Q�x)o���pB۬�s4
�ʲD��~����z�!�f�8��(f�w>~�e�F	�����'C^G��lC�:��¨���r�L�>����y,�n���ϙ���cGt?�j��i_��ȃZA�R�JZЗQn��\@kO��A�u��(��P�I� ����OH�i�[���IQ�ː?}C�x��	�B���v��ǽ�� ʉ�A�~(=7�Yy��0�e��Yځ�