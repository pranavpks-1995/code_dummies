<~D\����'f�!P�X��6��C�����A�QI���*Y���7ӥ��2	{(S����k����
2-��n�����ϱu�`rDk�kU��=v#�ӣ�Y���O~�[���߂�H:8����+&����M06��^�*����~��,�P��%$�gH|n�3_�cJ��3v�����$Q ��(g~���Ʉ�3��u@���͇I���2`��N@C�A<�\���/ڽ�c�I��"*�F9�e���"��`ץ���b�ul���9\h��+������|<n�͟�@�Ѕ�V%0;j�W����OtjC�4zQ�� Ѐ�f�E߻e{�����TDl�)$&'��|�]�;¨���i��,����	Ϟ�5�9͌��}v�p�8��2C���F�(9��>�5�Hkg�T	:
b��������TY	"$MJghƎ�ۀ�?}��Sfo�Cك���g���9n�̺2#U������
�g:/E�rg�ʙ���pskf��H�2��+�*{������$�|�9Z��Yk�%�[$����T�>t�TE�[ �a[]�4�c�ܿ/ CO�-�1҂=��N��.�������4`��p	^bY��P�n�l܄)�����Ƒ q�}����-+;�y0A��[sl�D7�4��#}k��Ǩ�<��g��N;�����6#�� �S�8k��b�-f��77e�Q���0c���l� ��zq�Q�t0�\z(���܀�Ƶ�x��"s_^�ݠV�+Q�$�aϫU����k�Gb
?�
��8�Zk���QFF�@�nh���xd_n��`Ȏ����
$W�U4Ζ�B8�g�2 �^���!��G$8}&�GD⼸�9{�����/�̾7�,���O�C`��v/�-Y��j�ѪD$�5j|�`�^v#�Qߏ9����S^�ė���v铄��z�� �;՛e��������0��ܞ����N��נ5�����:���f� z=,���M�U �X����TbxO�b��j�ݴ�av��s惙�a�>{E�T<	�
����4~"�Z|���R���S���W�W�AV�	  N ����,taԖ(f	R$�#�'�z��m�n�L� #s2@1��~�7l�����}�MRS��m`���Ɍg�P�ֵ��x�WD��%pJ���c���ˮG>�qx�h�q�.X5Y���$�ӆu��v3@e[�\����ua`���d�i�O�"�䃃\[�'ӥ^S�E�"<-T�D5B��>:��T��x^�>.�5e�kܨ(�s@t�q�\ϟt��Zp���e�`���Df�E���'�O�#��J]���W��3Q�`lh1�M��T�Ru�8h��4-��t¾��w��׹X���>�=���!��B	K�1f��\���eX0pPo�]�5�`�A|�\   t ��-W����,D�fʎ*:��j�_ˏ�-�V	�(r���"{�a��+U���i���wU��ߑGH��
���˷Cd�m,L�f԰����8��F1�<��M��uJ�8�e�����P?yxʐj\��=����=�u�7��G�5�����. 7�,�;���-ȥ�;�Շ	-�5/���Ǟ�K"���q+��E4�@㵠�aO2,~��;��aő�Ɋ�6��t�jX�Y�H�]Jv��|9퉁�d�G\,���%��Ƅ�r�����5���F�
w����I�$;1%,���8;<�K7�o)sM�~���Vx{��N]l�[eo��ǻ6�{�-{��!�.���apv����E�=Ғ@	���%Χ�.f�Zp�R��-   ���UW�C���@n�5�DK	�m$Ǆ�6�-f���5\+)�ԙ�$PM�h"�9�(��N+�9��'tt<N�A�1[j[\5�|e��yK/���F�yMM��;�4������������ˣ�>�更 �#x�Ņl�GD�m�r�q:���t�'�����$t��r�h�����Ou��1��/�J:_��-���ۓ&b���kF7����;Jcx?�{�MT��rSG�����߮�&��YU\��B�k�&x��;�F�3��1<Xo7ܚ��, ҙ��-Ǧ_EA	_� �=��?qډy���[�SK�Zh.�We^��u��\����B߉q��;��;?�GtΪ����s��?�GLج�/��&f�N�x%Ȥ��f�	gݘ��_ޠ�۲c���$5�����"�LFT�_�7�=���d>�p�-;��?#K��Y��" �D�� J6�$ǝ�����˸��'{F�����H ѹS�&�bwW�,��C��NJ=�h_	X���t�����BTfo(�W�$�G�^"��L��^�uֺx�݌1�zr�a�r1��^��eV���)&����#�>���^���,V��-�BX�g�����|������ bmt�$���-8�'V�U0�Ä�IX�K�1[��B���d�>�.X#Co[j"�h�bqB	��f��LgEu�dw����P��l���yβ2f���0$��P�a�ٲ`��4 �V�k�n.���%�1V�;JA�?��X��|Qo�J�!�P�_N�y����L�d�$������$+��]�6�32��w���&x���ZV���&��y����ԌG �@�V���Q�U���aI�M�>�[!6.wPȢUX� �k��N3"��f�A�^ݬ�f�L��� |���}ʅ��L��"SY\j�Gb4a?�ʲ��xf�d����i��>d��5������o�bf9�����y�9Y�<}�F� �A��}�i�*�8�6��`0�[B�M:�Jb4C'�(I��|sS��蚮>�W=�����ܔ��uV��}�7/�]c0���ŭ
�2�B�?3Ր��Fwu��I%6�lLl�ˈ�!(Uo�L�M�0ѹG��l�}�NΪ�Z�i����&#[�^ǆҔ�du�j֤�N<�)��� V��$�neKO�����Q"��
Z�+`� �1i;{+� )��	�������OL:�����-ZǅY��:�;���Wy�.����Xͪ��߱�CM��HG����f����T86@�в-jH��abgj�+���؅)��iT:�9j$��^�I�fhK��I4���o�k���%V��jn��ex�;�pT�9���TT�bp���?}�����SF��3U)+y\^ucM����5����>E���=���#!$P���*�\u��� 0�4����dDT����1��9> 6��
wi��k����H3�B��#��<l�|o�O��W̹���ڣĩ�+�(��;5N__�d�w���h���3:[&���CU�v�w"wX�����n`0Csj��y�G���/Z:Y�N�λ8����5�7�f։{��G7a�O���Q�E�~l������2�����vM
sd�����(�qf�D<�G�O�
�����]<b��K˫���N��|��1xX19���;����� hw<>��[�`_�W�����QO�N~����ݬ̀nR_��W���r[�*�T�;��bip�.����Ω��~�	��B����qzݯ���=∯̩�?�.����?UZ���\�����ǈ'=Q�@�I/��%���3�-[a��vF6����������V�p���5ʀ�aIuZ�2��K>�jn� biOK!�[?A0�%Y�t��/k@�Y;'�_�ɳ�9��%���[�,�������>�|�%�񲪼�@^����e�eqi�;�dr�FYR���2;���lx������3�':z�� y[\�_"��>8Tq����y;�#"R-o(Q[Υ��a����*���xP�:|�p��RMw� .�F�ny�-zY�c����gcG��eg�Q(�E��0JZƘ�U��툩�hބڒo�1h5��j3^%�M�y4͚Z�Le3F���45R6��wI�T�w�&8��*��ϐ�S�b>J\"��R�U�^��\���Fa�b�Vr&�(3�!���YIY���8�x�����3��=[����B�=���Mf�arF=(�.(7�v_Q�?怠V�����k^U11�K䯔|��wĔ��\����e��|!pG�{�N���t�α��� W�zFo��>���F�
j�(��}Y8�*��-7N.���)j��[�"Py;뿩����)��D>0��B��#�Tu���E��.���dK�E�G��눆$b�� l�!&����"n��c�����]B��m� Ლy�t�9�h�L�*�#va���^b�-�kz�M���)o�,�]/Z�������Ʀ��xs�/�����c���Ώ)Xk`�vՄ7����1�t��+�X˳[-�h�q/_e�hN��VF�A��Tv:{��[�J�75GI.׷�.�b�[/k��Y=[��}���j>���v71Pj ]4��jEܔ�p'�Σc�'~� �1�&���a��'�f�C wC��cG� ٭q"��H�S4��I���b'M.W3y0�N���i�tu�|b��x �θϝ����?��V�Q��JΛ�ʓt#�w����1�rd��p�!��Ei�n$�ˏ^�:f{�y�8Q~�7�=��v�o�bF�SKX��n>	�����Bq��0��c�M^�����������4D!�[��[��������Ʌ�\�ѡ^��ZuZ�L�xoM�y.F��+��KWO3�'Kt�l�Bsv� [K"]�c�g �mz-�w�k�U2����m���Kp�m���{���1�Ñ8�ऋ�$g���W��v�"������ˋ����=���f�=����Y�$F��D�r賔��Br�a1ã{7�#�q�	���[�ӣ^ j��&�JG�V�#z�ڴ�\�U���m��VE���g1 b�	 �x.�4w	��ON��]�'$�>�~:�b,[��B)�ԓGУ�q(?�T�r��?Qb&#o��颺���T�b����y���ª�bl�	5
!O3k��Fn��ٜ[,��,O��.�J���*��@ܹ�ۙZ9��^�z~���}�(�OY��6A9�� �mbE�E�6�py�"`3�`�]�>%;6��5�\�?�^)ߋ�����8�v	��j�	��Fޢ��-��L|T�܄�n���-��e͌��@5p-�
�W�yBF�����"w޷�l]��w�AWW<�9S�ASHR
��d��Mh ���U��̧.�+�^�	�z����i�k�*���CW%?�^��]�Ń _�W8��:od[��a�
Q��ֆ�J�ʴ�d� j��l�G��3s��k�b�1�����Tͅ�_�~��g�h��\�2�8���=�B�M�NU��u��!}=u�&�ՙ�(�Zf���}����2���Q��B9�G+<4��)�c���?W���c!�d�;.���T	���q4e�#�������mg����4�YX~+s�f�$��^����9�*�����q�s�o�Qu���kP���-+���0����a�rz�`���[N�`��VH� imP�~�����/OYîB�eg�N˴s����ը���O��T)���_�e��x�H9��fԯn�,�5��=i�]�d×��g]k�N��M����i Sh%���lv���涀MTm@G��fiOQכ�Fv�
��ߡ��7�ZN�s�ˢ�GHIj�3�ND?�5�FX�`s�[8��&�Nn� �^)�u;���V�i��\�4`_���p��IX��� U#��S8}�W��'��e]��֩ϔ��O�1���Bu�I�Y�V��3z����ӼX�ʂ
&���gUN�=R����"A�K@��qe[�e1^���]8V������&1�9wrZ�}�	2_D	�Y�!Q����e�W^,�T>o:.E�j²k(��+s���ù ݐ����6�p�2�¶yx�X�B��u�jȂ"l������ǘ��/���.NB/M*~�,�W���#�9��i3T�2���*�T�a%w ̀���'+r�4��k��M�.�c�q��������⺣���Y{�bӒE"��`�#�	�S�g�EU�鵸�lh��h9����ϭ�DF��^�o?73o�3�jg�k�ب���jJ�� �r�tB����^��d ���F�Q=�ike�K��oq�j"��Eh�&� �ԑ��(�{8Y���2D�R8��t������p�L�� ��qw�{M�¹�߈����`�"��K�<.&#�p	!0���Ap�np�����W1j��]s-	�Y`����n܄s�@�1Og�9�\�<ل��c����I�MZc�nx���+��O�Z��?�G��~��k��3��Ņ��`�?#Fq�嫞�-��+�<�O�W�o~���(�F;�Z�A���X��G����!��1�g�����V����^]�����4O�z{m������8kF���~9���?F��A�Wf��@4�d=�H:<S���=�����h|�z���v,�}u�Oj���!^w�Cإ'	L�֣G��  ��B%RW�c��*�)P�I��+� �k�j�����M}��@y����{d�tg&�b r�ȓ	o��Ѓ��u��3G\�Mm{����irc=~쌣f,�#L�Z~�"�_����,h=�h:7΀F����>����[�mO�b��8M-J��a;��"Q����%�,�=3,v�\q\�!R/s���%�S3��Dķ���i� ��Ǘ3����^�-�]W�%�a���7���YlNn��V����c�`LV�3�����H�;�ۑ�cC�/��"m;�<6q����]j)=�`7j��&ݕA�����|�#�l�=p>4��?w㬠����䜫�r��M�� z�d����ݫ��CF߀p��HAe�W�U%T29�'���o�X�W��ȋ�ϯr�v��t�@���������Y]��Ɏ�`�4���^��Jx#�X3hWB��^.Ag�>�Y��-�TyW�5����h&�{��.������8yqD��G~�qc����{~��iN�'�S)�>�E�M��Uj8�)�����6nZ��Z�"��>O~���Pဳ���j%Xs���pq�I5T���Ɖ!�6*����g��>^K��UmP���x��FΨ%�jҞR��HoG��J'����&�]1to,|\�bN*�L�e���gن-ê��B���X<�҄ę�B�,ٳ��ēI�9��GV<��!e�����i� �|B����D���H���u��P&h'V���>��^~]���vC�l�Ű�Al��	��c�e���:�d����y9���):V�kC�/��w$����a@����7�G1�Ii��)"e�z�C#��!������2���|�ޠ������n;2�J�J�)�+������h����E�S�߲Ou����%�������=)N�7�0%C�%��7z��� ������3�Nӄ�jVLuU��Xt'!.7����bFt*��_ַa"��P#4.��g}�@�5B����x��O��o���x�<S�β�MQ�Se�/eu��y׀m4�����f��������I�1e4�O;��Q}��O������ ��`i��jfq֝��&�	���RƝ;�~�C�.���f�,&s��hU�%UH�U��D�VոD`�`�4B
=!/6A> ;���o�F��l�5B,��kP�I%�֏�4u@,_�~R|^
�'�����bP}��u��'͡$R�C[�̨!�(-'�"�y�/D�Ɨ����-�bY�ݢ���+:�����kmK��A:
a�"�%�iY�N����C�&�2��s[q�C��jDH��&3�]m�׊S7�%��F0�J��W"]@�6+-a.OG���A��$}k��N�	�{�^���5D�ON#\���#+H>���e�-�טj��0�CY���k�"K5� q���%��ZE�m˟7���W���дl"DSN\����`H2��E�HĆ��$� }�$WVu�s���[N���9����D�C9Ma;ƚ��/�rW�U�[��P�{Y�� pƍ��2s�U���'b��Q�c�xϠ�{UF�i���Y�U'د����=¨�k�p�Q���Y*)he(�K���9
bYJ6�,h�w�I���Qc�S~VXr���ڕ����{�(�9�@��������D$��}g��Z�8����|4�>����ab�s߰��3�:%*�5�ho'��Ψ\º����sԫi�ڣC���  ~ �&���,t`�Ƥy�������M| �u瀇�V����b��:�'u�=q,%e����"�^"�4/zu��4���1M_��so-�MF96���\
���}QZ��V�K���v�\��y����8M�9�˔�Q�#j2ùLe�J�S��D�{X0�U�?)H^ 1�YM0��et��'�.Dd�?Y�