�<���q2���l\�T�xe����(�[v�$�W��/Kj��]ؾ��e��J�����eS�U��x�M8Y�fJŖ"�rE-oA�xt����q�V�#��Bw/;ZRxi������ pLe�g;j鋷��U��uJ3	Ѐ~u�0;ͳ����\C�r�V������ t�]]{���<���m�_��yi �g�B(7�������J�m�d� �G�ȷږHl@�T$� ��H�ҷ������Ԗ��Ҁ���h��湇���0s)��i=���TM�߂�� �,�`���y|0��K�*��OpH���<�q?���Rީ��gB�b��>>W��',>\��c��_=��&����M���h�z��a�~�I�J2�CKyѶ~���"�:��{�a�V���x������T��(,�0�Z*p�n�H�}m�ɻ�+7��.�6��Q,���f:�W{a�Vn���W���ȷ?����7>��Eh悛���Oj`�ew
|oaf�y2\���cy]EVhɨK�����m^&Lp�Ϝ��h�3�@{�K��}#���
�<4���Ki�8YzӺ�ẉ��FſVvf/�H$Y�Q��%�[GUĈCb*�Z_Z(����Y�O�)�I6��'��k�6�	��"���14�bd@����9��Yf:��cf,�O=y�۬��#Ó'��M��Qb*�������d.7�3��WHR�@�D?�M.]}��9-�=9^�3���z���;��FV�ުIg� .�bK�<&9	=T�-��u��Ș2�&�c#�`Y/��.���2���Y)�O��5}�q��'���� ���QF~��8�A�����������{�@/ʃɼuaՖ��T����a��)<BAh������� ��j�V��x:%�E�˗®��;k��(��0��{F)Ye��y�:�u�:��&�ˮ|��D�S���V&bR)���TZ���4��*�ɫ�o�
�z�R��q�>}	���\{�[vm�Ø�'̅�#ߦ��ϦV~�f�Wmw�}�sӉEKx�Oj	�ƈ����Y�l�@�)��o�o��s�%,���Q�r���
k����D��V(�,�k�u4�?·�|��lg�*���&���S��Z�kO�tʲ2�Oxߓ�T"��a��(g9�JR˂�����+Mg P���¡6�Ϻ�i�K<u�,m���<��g^�չ���k�9�Mp^��iul*������&�,�³r�mn%�IE�.�,�Ar�H���~�1_� o?�교쩀z�@�^f���/�P$1�z��-q 2��
�=�#�x���L���hT��Aŗ�Mev(��
���S�X/�X`ơ���V��ix{��d�Z�y���db#���|գI���kh
�. �X��+%^�
���پ���1�&�:�;��%�s@m�3��t�38�ۇ%�A�e6X\v��@	�g)��i:��_�E��G�ꟺ˽0�����چa|0ۣ�h�P�n��:�p�,�+�xIRހ�T�l��:�z�v�K,�ewX���0�R�hk7�j��J�܎d����l��uxOG��e�^���n6�(��U~��?�n/�:�W4���ǫA������EZ��.�u9�����th
 ��'Ah����#p�~�M�*MÚM���ͳ�6�k����w6�Ω��W���aP���W��:�ɣ��:�!�C��(cc��`#%ԙb�7�ڂ�D�~o���������O-$q�gM��EF���M_t8����s�Q� �ɋv�4q����v-jS��"��v����x�~kq����;�CG;�B���Q��K�I�ATyW�Ȓ��0�$9g�y���3k�L=���K�$�]�?r���%�[�xU�������:���B?����rR�&K}>����w�2���?T~�©ph���cw����CjZ{c��ң����U�-��ɏ�$/��SȬ%�Q}��&�$Y&��)�3���ͫ���ѽcO�{�l��A���o� ��ɀïݓMT�3Sq>�+-�G�o��Q)-VY�m���,�M���0E'����]N{�E�� ,8�������My��R>��u1�Lo����XR��N����@�KB�}ؘ��}�YP��Ï]��4�Ƶo&ic@&eb��*J���6II�d4M�Z7�D@�a� 7��b�ٝ��˴AMQ���v�'ݩ�4��9w���;Uz)D���t1BoT�g��j��_ؿ�*�
l<苖�\�����T? �B����0�&a�g�W\�M��T�a�f$�����/�]Cu�B�=�ʝ���w��L���Tte{~XN}�� k:�	(F}
m��R��.�㓆��V��8��P�{�3�!��fP� 	)��`�dV���p%8]��4�HW4�p�c9x�uo)�=�[���\�7V���C�n6?�}�-2���콀YC>�����]i�h}a��l[V��3�����Z�;�)���+૰S�!T0����F,naM�z�:�s!1ᗤ~,m8��Fđ6׵��ta���n|�"j�:���vS�9��iK��ur��NM�^H����5�9%�X���
�*�Q���(�Bu<:�9���x����V<�3�닮 ����cv�"]�}�O
�� E_�c�n���k54&ٿ��4\�����U=6,O�z��k�w�ȇ�g^��&Ĵ��|{(