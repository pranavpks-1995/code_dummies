'h۹���#��n8 ��{.��g"������\��~�\�;���I(����e��Ǚo�+�J�ȴ-�7N����:��4� ^��_3�Y��A���T\������j������E�\�:������î�q1/qJ���-�9fҞ�5���x����E$���H������/���*�&�*�H_U����!̏'����Lp�2��ϕp� 1�U�,����\�A�����x�_�?���,��욊�x�S�3 �L����E������R���s�� "ZO�.��!5$�j����B>:�	HKQ��{��7��of
E�vQ8J�mH�֔{��7���A�/L���G��3ql`5L:���xh�ՠ�V��cHY��J3�COqW f|��2$�Q�0�ԭ �k><�M轞�$?U�>��EP�r4p���,^��/�Z���N����1���2�;3%���V��π�ք����������HO���o��uU'PiA�ZBU����Z�� ���Գ*�y�!�����4���c�^��^���q;�U�)䉮�|d���6}>o�\A���c�dQ���̧������e�p��x�X撵�J�#蚇�V*�X����7n���?F���<�X���BK�K��zRjƝ���e�ܪ|ړ�lc?xDG�$>����4�Sx��#7��_��<�����#�x�=XV#f�*���P���Y���kiu���2 TsR�����G&5�`ʴ�B]����E#�PRy�3.���%>pNy7�_���J��������i���	ĥ̼����;B�{W9ԸrтSX?ց�e|�t�GRL$�/���a���]��-y�6�!
r���F�N��.���tcx��*��f�z�I��z �o�m��b��/�d���\��`"�cȆ��!C�F"0U�uǰ�hj���������y�d�x�~�����K�Y�}��-��x�9�Z>ӥq�s�6��KX-��`�Å5�9o7K#S�+Ub�7�*9/����#L��g�i����L�7tJ�3D`L���];z��C��I*�4�*�S���{3��	�"�L�}ز�NL�ӻ�L�1��'~K��LX�pE��v� �t�EVW�