P:t�=j��ڹ���&�\ۚ�]�~& ߊ��'k@6m혍ﲙ_�<�D�})�W	���L�����]K�7ІV���8�=��3���뉨��'"S����ܨ����䭁��*�S�8np��Wa۽C�V3r�o��5�R��(���SNM���L�Z9�ڻ[P��R���dI�ꠛ�KS���J����ى�Φ���ʭq5�Q����D��	�ż��xw3~��721=\���[�aH�lʳ���CS��kA�+<au>S$Ű���ۡ�-u�f��W[4��A�Yؾg�H]��H�x0!z?P �w3�J]����4v��[j@V��8�>��x�G陔�u%D���:\E�,���-��#�rR@8�Hֲ�8c���^.����W���y/8����n%S�̡ɖ���_�[�D̈́nq��/@@u^��^�����zw�(��:��u�]����A�bV �ea��F�`o'���},i6Tp2|߹��0��K��5 [<�W�e��l�-�.��3���2�!TE'(|�͉��~BP����v3̞~� 6�1{h�-,6]`��� &��j�/�!J�V�%"]���J�ݼ���H�r�5�S6a=N0z���/�d)\˱Q
w��r��]ԡ8 �-�ڠ���U!Re�^���-�ƻ@�g��s1�`HB�)t�� �om�`j��ߏh0I�I/K���:;"Ӏ�ED�L����Ȥ��!�	ƃ��2;�%`���][vd�KP�����cB�Ar���g5Ft�J����5$�����?�I�Gv҄�61�V�usf�鸯�@۞f��n�W�Ï�xpSÇ�s!9��:��K���v,�w��F�	 '��x�&I�H�Q6V�����H�  �!�����!���	���S A���O��)���v�;uU�d�x�"樸�%9�Ϭ�F���c2�.����X��CD��@��9k����a !Q���\��룯�R \�.�!�5�(�'�SjۻHB3�/\��(4!��=H���H�"��W@�,!l�����#R�jx���8��A-4�D�, �:��uߥ�� N1�Y���
)Gs�]E�Ctf��~��|lk̀=�mħ\�4�^�L���!o��d?�����y�γ�a�H�~�p.f��B�}��R:v�!X����=|h0 �!������*��! ���@`dߡ�}b#ѿaP"����
c���i4��4�ޞ�H�>�땷��θ
�_W���f��H����i5���(��vi;�(goӟ��l븣�1�`�6~����j*���=��6
��D)
!�E�5R���uf/�� 'L����9�M�F+�yV�A2�� 0   0 !��Ąp��*q2F��A�^Hm��D�[E��89jC�D��ąB���c�R��B(3���J/<�	��� �ᙞ֯�{<X�Թ�����g�@C�b�ǟ|~�r�-�&�> -��"&�Iw��NI/�)�k}�������w;��|�0      p!��#���PC	H �E��`�]r��RF��"������U�)Y|=`	3��V2�*��>?U��TЮ����@cu�CGKF@��fS^�!Ean~�VY>㷫�[�J���"|��~�\ �P��-�9u��J��t���^��rV�`     8!�
��!���4�X� �  �R�i��\* �'��E3 ���9��3/��0j�� ��7ޓ׭�_�<��폎�s�2��{�i��������8 �� �E��  ��)���$����奔�����;.���#L0     ��!�+��B��H2D !j��Z�l˞ ���$��[�:A���M�D�Y�]�T4�M]�,��Y�{���5�T�u�K���vx�8��
P
��B�(�k��4���ȷ�v
��z���A���k�G_O8��%��>u�W.{x&�cw���V�Qtr�    �be�y   "]��UW�C���)W�J��`S0����1�g�����bN��mQ���n:'�1l������b盅g��
���G*�us�jk�g�"��F���L
�f`�ZmzS���5���ߒ��_���DL7�y� u�f]Jli������G16����D��;xA�lj��Ŗn|lZ&��N-�L�7-Wű�7�����!�a�X�-bfS�+�N�5�2F?��(!����-m�p�dw1��k#��� �td��7�g�x�[����WE\�2�Fř�O��2�ʜV�%�$�Q�	pl��0|�h��]>H~�F�[lH��`UWAhAN�n���Y����\�{�F� �0�١���1_�O֓��.���C�SE��S��&2�B��ǭ��J�i6��d�}�zO�c*�B��K;?��jQ�Y\�x�[�p�on��o.�8&c\`!�T��������:�!C��Q{`�ͫ����"�[lY�Q�G�YX8��d��?�+4~��8<���@7��F�tѧ�n�I|��6����wh��l+_�z�7j��36G����(�2߼L=�������?|��f�4�I	0�-S����;�Q�*��"/�?<��=D��?��O������M��83��B�]�<�*c/Җ:� �d	#�������|Mo�e�i�/ĭj�ג����T�h,
�^q(�P:W��W�����GWq#��0�U\��V!���:u�ex��Rc����3}�8�R���T.C��3o'`��cHԴ�{RCoZ�f��+n,��j�A�)!��5�N�\��8��  /�"ln���I��h1*X>�a�ǰ}2��REs<�b�+Jg��5�P�t�/��� aM*PD���[����򀹁ɡ����pW#�'�<�h�9� Ih�z�����t���2ⲵ��h,7B��ջ�����y-��з�j���5(��8�5r����%a��Pi��S[�Rog�0hf�d\D�#T�*���B�y~�|�qw�=��ڙs4��àly@x|��#��2�g&c�4��{�K��J���P&��S�cXɱr��^E�-����?GRV�؏HM��b:M)4�U~΋��\	��IH[g��`�{+�(s��{��BFOO�����s���I}h7� ��)x���S�Z��R�K<������_��q��a�mzC�����qYE��"���)��}�,`�i��������ŷ1Q{����C.�L'����[�:��=���=1Z�JSM���,������? �~	���Tdѩ�ɛ{F�����u�!�V�{
������f�2���ܫ�/CqO���OVz��S�6b'Ic��o��%�(�G�����Y��;�=$���w���ޘ�o~��obB��0x΂Ӣ���t:0F�$t4��Ȣ��;��j�X��dd�<ײq	���c�Hd������	y���e�Nծ�R#�>^��f�r��^�_,� ��i��Rn�ٵPԃ�̓(P��2vP�H��|���D"������d���C��@�D{�w��恠@�ׯ��S�%ub����޹���@���pu�D������1O�<4�Y����\�-K~d_$Ip���b�3���Kd;���(;�6��
r#B�x\)�Ɛ�:�B��i��1:�3؋�	�b�G��H,>`	�0�#"j;�k$�����E��J�/v2�UB5��'�A r�4�CB�{y���C2n�����A=T�C�dޜ�YY�E�� �t�/m�xHG���3a�=���5R�=�Z<ܤ��J�G������	M��!�%����9���C������{�2N:��HQ\3n� ב|!
&���eP}���cf|;5t9�Tv� 2E����К�h.'��|�q#�|����b7�mZ��Vr�oA�J1C���t��U�Uo�Jk_�=@�L$o��D�}Z&!�vDj-��f��E.���ˤ4\ &��J�h��M�X��LQsp5ۅA" WsF��D� h�Sʾ�_U���� ��K�s?km���:�Z��H�('��׼Ȝ��X*J���!"������yaQ�j��Ҍ2pXo����^�:�]?���}����W_���̸���L�V��BVa�i ҃t"7���㻴���y&r:Fx�Ud�;�Ύ�u����ڿTG}-Z|�a��R��� Mf�GK]ǃ��K��w�y��)nj���n�ޘݒ=|�� C4D��z^Z�^{f���"�ΓI9U������`Vً��xB�"�U�b�������G�$h��+�ZN�p���Ab7�A�9m�.^�јHD/�FV�/�d+m�qP�������Q����I��/�+��&�Q��e�ﴮ������YZ�PX������%�א$S�@UE\�%�>�>'>���Dx���gN���;����uy�h����y�a{|3�Y��.����0��XC�����5��2	Q97�d
��i�Er0�lo��(o�B�!^H*j��Ԗ��D�<j��ʲ�� �J8B�a��pK�.�8}u�Ϸ�l��ٝB���`c�$�q��Pژ3EA�h{4�u������Ds�� T�OZrr1��r��}s����QO�fS�]R�!n8+>盭�a��U(������e�g��6��(��a�L�ћ��Lě�Ò�l�����#�ר�Fpƿ|�݈�e�$l"�/��ƖF��xC�w���2{�K�7�j��(z�P�N���������S��V1�z>ER�q�n��+YgRl` �/������gd=��d�_�o�l�*�Zl�R6�y��5�Pyr��1��h�i
'����d����t�:���9vs��*��[���֥��'�~��~��Z��=��,v�r��=FŻt.ӄ��O^!׽��ga9!��pjk�N-M��W�n�H��FA�96(Wq;ҳ�R�c��4=��K�b�E��vl$��,C�!�ƞ��l4_���ȯ��YES�FQ��I\�J�c�f����w]��ƍ�0��d��c���9��n�78�eT�d�ĺΑ<�5�6��_8�aH�0�&!.�ԟ�S����F ֎�zl珈y��o�$�UY�'tb�/��~�J..���/��G�U��(��q����G���E����@\�j톆��T���A���=ɰ�I��cو�"ݻ���3�t{+pYU�5�~�����v��͚�yܱ�'�ed�<<�u����|��dL[5�2���,\�b?��|��x��=�2���Ŕ��Z<�9^>���`�@�yӜ;61����*й�i&���Ô���ݳ���Iz�� *�-��v���H���h\P�up��n��!+|
��Hi���ͭ��%�4Xk�r���~e0�XH�3�o[oa��V�H�,�zms���ړ�wӗ���F"��@�N?#ա������T�؃Mg������s�^Xy:g�5�Y�L�k��k��k