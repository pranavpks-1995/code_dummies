�4�05�o9i��Q5����Yf�̼���ib'���!PŘn�3?��*r��7t;��Ì���qf������\��<���7�l�!�C��D���D{��ؼ�6�ZS��xL�ЃFr�ջ"� Ū	gɂ��-������yJU3��l�.�3�AL}�x���<�/Ɂ�
t�ތ�	)�o���쏇�s-ׅ��[^�@#���H�@��6��Y�B ��;�T/�s��B�Q{�k�<��a�"v,����?g���Lv���,�v��u��R�ֶ"q%;���ؙ#	y���ۖe�P}���,*���o]��4�����Y(v|�yW�mCz�%�����z�í�l��6��.�J�h|ĳ=K��!AlД�q����#��%`�$4}̕J��bS�$�1��~���Q:s�z���<W��r����;<$�N�o�x���2Kz�F�Y���"��|�����OH�"��3!�h�4���J"�������碟�,�PM��s�d�5�����`�߲?.�����2/�o0]Zd<B��(��=k;�j=}O `�A�u�������6���Q��GY��Bg�Fqkj�a����vRi�ʚ�$�G�B�?yz����X�q��~����lJ[:�1����l�eG�Q�n�'�K'D�d娉5�pH�N�h+�{\��V?�7�� �Lq�/MJm$�WʷA��	=�����˵A�Fʢ@P܌[����S(s�UA��0�����Z1K�5Z�!�B�/g��-�H��wt#=0��K��E�m��wB8d�ڳ(ŻP���Y�ff*庫5U:�f7DKBQ,ݰ�[�ǚ.s�x5�IaoDi]x�(���FnMU��	=+���o��į�=�r�B�@�6A[ȤO�����Xbڇ���B΁�  � �&�U�#	��̴���|p��<�M�m��7���a?���hL�������f4�8������vh�L��ԓgt=ƻ���N�;z�(7ٲ2��%HlY+��Ɠ,�� ��y���S� ���׻�����er'�N�������Kg@�D�I.!����������{h��/,����Yf3L��x1Tsm�܊����p�������9�����ɹ_��u[�H�kl��4�h�K�]&����i��~�����&`�kw�܊�#򿆣_f��3�� �8M�=k����p�Li������mkOZk�m���h����ʿ����ұ����?ڌэy��ɨKL�G�Q1dc	���`ݫܹ�5��p}.k�JP���Dί��t���T����vzۄ'��e��(w�`m�D�@,L44��]�/1�5��0.<��%J��/�N�]���'��sK�a�p��d��O��a�J�w�r'�E0�8�-X�q��wX+Aԥ)�2µwɎ=��YM[�X�a���^�׆�z�a�m�9gG"�-"��lY�:�@{1{����D�s�s%����.��)^j� u��#<���,����C�9CX�}���FH�LЉ��ֲ3�K��Et����p�:4"P�j���JQ���[�h�/����K�~�d#��w�F�B���   � �F�u�#����𐐔���Yo:�8�V|�!��'~^>���I}��U<;�j�=�}���$�UW"Ȝ�.��8����2�a��fe��a���	t5�����+�	h���S�ZGyU[�c�Kf�^�p V'�J��Yʑ�1����A[e��\�����WC�Tf��e�d�M�U���!kR�-$pZѲ��g9mY��l*D�K톮�u��g�(4u���Ǡ�j�V�ыL#L�`G!x^�\�Jrt F�Sd�wn�_*7R�޶o5)`�����Ë8V�P�����g�"�֊��Y�N$�|����o*��?8Y�4H��V��w;�H+~��Z+fS.�������d�:<��c�ťQ.�N���������M��-ӈ��u�_��w�c�CԕS]FLA�,�t]�Y� T2v\i� �P�%K�g� s:��s�a��7l�r�L�O�0�����5�����-w4��dAWʜz/.8]�4��ba��sM4�̷�6�t���o��\Y���owy{�p�.��BĲǛH���b��%׷�F��f)�T�g�Fr���s���Y�3��-�<�#��G�efF_�56͚�����<�
B�xx7Yg����<�M�d"Z\/q���G�zd��t�`Od�W��o*�@�C��}'���$yȱ��;l{�6x3j-�(�z�@�-�>0�b&�����O,�z�)���gJd�o��`c�G��	7[�7�䈴�(�?���H����A��   � ��-����Ո���(�� :���$BM�Sz5I/o�J>��]�fO��j@L�L�ϝ9�6|:��/yy?����u��'��N���P9��VR3���V�"nrlk�8�]���@��j�0au�)-WI,]�G-���1�eV�
l�%�xF�,��^�2��%��]V����.����}۰M��tcˤ'��#.������P�G�ʄh|�0��~�sDSG��G���}����z#��WC���:U�2�^{���(�U)8D�s��'��S<Z�l%��*��������v������2u1a3Y�lb,澯�K�2�m`��h"�.��$�
�a�k�����J0Ϳ<ɜ�|A�'�X���m�u����8�v�!w�K����)<�+�C�s�WR��ހk��]kP������ Okay.���Mȁ�   �Ո�U��C����Ʃ��B�:^ ���n���������j�1���@Y3��!�"{�D$��p�~�s�P�U��7U&v�3QU�J�#v���6(�  `=���{���oW"N���º��,O�e�� �Cg5R�6�t ���o �����~���#bnN�%��N�=�&b�>�Q#�B�s^�*�p)Ԗ����U�!D���mF�XX��T^���]\d|є/(ft�^��hX:�b�K{i��M]7�W����6�su3D�ѝ�M����	K���j+d��}�H���9g���:.-
٢�ԭ?L���]Ë?�w�?�D`��U-@�bB�����G�:��p� �}�!���V��C�˵�H�\������G�1�����	�=�E	������Ip��֖��D+�/��+j�J/��P��_'��CX8���[�v'�8��XYN��UG�$��L|��l�as
�Ă�8B�G�j��x�B3���z���m�F3b�9�.i�������<�)"���T/Q���~��d�*�7�э�H�ɯ�ቖ_�\)8O���ե��GtԜ�V��>���)��rh:�ɮ\�6}�8-�{��R*VgD|o�б���\����M#^�ͳzȇ�.�W_�~&��U��k�Nf��s��؃�kQu�B�#*�5�O&ZN(Qj�k�f�p��p%�t����uӓ��-��y������E؎T�+p�,
�k�07{�7���P�]���3U�{�L�.y�h�AƳs��mo�/qB?���-�����������ܑ����ɷ��7y��g^e'RZ m��?�*	.�*��8_�L��	
`�E�M��N��c�b���Έ�y��ܮ���E��zx�2����'�e�o��%�9��iۤ<͹5r�h㚴m�j�V�x&����*+s8]��#C