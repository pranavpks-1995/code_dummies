܎p���mkO��ϴ�4��E�w�c�)J���m#�!#C<h�g��X#��bU����W��crz�
��W(S�P�\�N4�O{	ˀ�w��
��r��S�>��ʘ��p�*��q���{k��oΤlT�����t`p@���]x"�|�ò"��������qN$���|�i���R�yS-ȝ�Q�2�	����~G�4u"\��v6���T6�_�/�S8�*�W��vu��so ®�b��D�����!��S���Y*���U|iF�F#��x�J���Ӯ��^za�iȫ��E�4�����O�R+L����B�pr�lAj��F�(j��}񺧤��T�R�#��՟�����<�����1�]�.�?�M���k�4S�v�;?�ՐՓ���6N��X,�T�C��}"47sL>�Z�����K8�0�	cDI���~�h*�RF��[�@��V���B��A�Q��	����L�ņ3zO�F7�GP@��8.I�eݱ1��)���K�R5��GbҼ�~��P�˸=���s�����ۥ¥�J����2.i;����,lg9�c|Q�uңB���  � ��U�"u�T�|D<�$n����W�V8�=fL�RF#�F_�T�($�ա�N^�t���j ��I��O���~������G��(�hE��n4!�+?q��10;���H�-ˀ����-67��~���t�Hx`��6�8��@�����]��Ô�%�B-��幵o�_���l�A����s�~ZM�yv�BZ��[�X��O���J���}�t�
"U����Tg���v̄2"f��%@Ey���0@A�{�����n��S�"�8�T�)4�{QJ��*�k���l3�������T��*�\<��'A�d��\B�J�O�&�h)o)�]� ��fۺ5>#�R�%�7#�t�H���4�0.�?�)���p�ĵ�v��MT���S�����?�ư���{���xKb##m3���_�-�����Pw�d��V���0~N�+��"�K ۠�� �z���w��PD�V'���f�t�Cg���ޡ��χwX� ��x��䬿#�
Ɵ�ĕYe����(�ѹr��?�y���8Pj��%~4�!�3���-c��EB��*5b�~��b���t:�X��Y\%�C0rw�M�ѹ69��]o~��+d0*��1$�-[V�[�31�a�+�#�B���   � ���u�#P�x�p,$X�z徚$kH��s��'�}�T'��0"t\�^��,�P�^��G� ��������Y�ܮ�A��X�y�>� �>��Hl�H��d��.ː��L���6R~~DヿYht��C1�1>O{�u��[�Difq���csޘ�Y|%}�"�y�~�$�4��C���Sǐ�Ϝc%u2�f1iRΏ'�ն��I�㔷8q5 �ݬu>��M���� �"���t@�qӸ� H�C䜿U炕w�<�@�/١�.]L���^�A��!�������P�W�mR��y�d��Ϲ�ɒ�1)�%�!��!/�E���q+�)a@ � .�B{J� #�H��t[Ӈ��$p����+���T�b:ڳ#^�>˜������)z�

{q�J1\�Aq�n����4^��f�e �D���9���ІR���M�ݙ�+�5��^��)��`ԛ�[�S�ng�\��`�ayM@��}�X_2�b��#��w�h��e��E(/#���x���J��Z�?Y�~�'�T@�p2����0�0�j2���w�b�S&�� ��@���-Q��Hu��I%�h�a���2�w�@O�v���w.�<��,"�Wg��Z*-��.
+�v�=@xv�HI�ЃC!�p;�S��\p$����G `I�,��x��A��B   � �-����琊��"�J^��L������ݜ!���+��g|-1ޠ�9)"��1~fJ��z'��|qb��q��bw��o��m�|�#"��.>%{7H���ss����iE\K�S7�B�dZ24^OA�c��ڜZ�[�Q2t��I�ԗ<�|{�T2��ƽ�L��g6�2*��G�T�uK�߳�]��\��$�?2���u�K+cn$956ln�	�ޓ�-��8�F�ߡռ���m�ۊ�"M���딞5S�"X�<�-�Q�Vz�)����G3�A��宝@U�1+7�^.��W�$�ƛ֘e�v,
���`�`�M���AN���m��T��^$,�͋&hv�ʱKᚱ��w�\�Rz0`d���2(4�-�2w;05��؏��hkz=,[�E&;@o��綉's�/?]�:������J&.�7؈2�,P?����.
/y-ñ�n�3��W�wӇ)qo�f���*�h��e�R����4��R��   zӨ�U��D:0T�X�����"�jc:0��.bX;$-���Cq:m��`BIB��9_;�V[�X�'%76s2���0h>H�C�'��z��V/ �������	��`nv�)�>�i�Jm��`\j�c�VN��jo<;�{�@���"�<{���3"׀XRM�Z^�:9�q~�,��<�%�{���MT|��[9S��DhM�[�}� ��C<�%�yo+##�i/���]�e���_�>���^�戝+;kվU0jI�kU�.W	~� b��Wol_h$9?`�|��#��#]��X�z�:�2��w�Q/�.���ZN�/~�)w��*�N�&�]�b��L?�)��a_):5����֤U��ь%��XjX�ۧ �ՅN�+�bGr�0��r��T�<��]_X«�ൌ�w-�� ���%"<�9*f��%�wL�Շ0�J����O��>�n����;�l��F�zqk:�1��aĆ_j�Q���/m�n3����P�oD�M%obQl��V�Ӹ�坟�1�ē)Dd����?@pX+3~X��S�	e���7P�,P�=!ؘN!���eI�'��'c׳f���H8zP uUxM|�~��[no��%'�K��pZ�Pf�^�AJ�촃 �c�K� KmR�.�s�YVΔ�W�:�G��rt��W�ۦ��������aS&C�\K<�����{����!��`�"��R���Ҡ(ͫ �_�/gh�3(�v/�t����EH��PH��[M�W]��9�F�1��h�k���ͫ���Ί�75�j�7p(@Ei]A\&a��^�v���� l�P6._0���f^�7˩�9�	9C�%j��h�}�3�Y��ٽ�4	J1�/�6��0'���'D��I��7�mo��^v{�6��{f����$��7����K):@��a��Ը���c��km�blQ��Ȕ��6�lW����%����83�x)�8E�V�$�@�J �4�J	��e���4c�$�D��eH���a3K����?-��3t9����˯
&��K�c�ɔ��m�9�1��:��a_�/~������<�g ~��t\�8z��Q�15�ˇjL�'�MX��n��u[�%�Uȍ�:�j�I�=�@��W�V���ݨu��ߙ�����Z��r�6�,u+Cdl���I��݌H6?�uЂ�X�Db����O�]s�0��Ww��p��2sw��.�ҘZ����_Vz$�g\ �yt����dUn��>=����|iC�B	���y̘�Z�W��zt9��y �ǀ�-�׳�1����!�($����܊��.�C��J.%���y�32	4%g��F�$*�.0�����ut\�OB�<0�Mo�qF�v�T�V�S��$��D�o��5��L>�6�<=X��W��X�у{EF�����'NjӖM�uf�jo���@�Sx��
�/&��翛a�ʹ��{�R��|�C��J5��nƷ9RfQ�nߦ�	u�a�K^ksFg�����]�x*����.�fq�`���T 5�x��X8�$%6FM���Df���A �#/�J�)�G�j	F�L�kB��:Qv�����s����f�Mx0'=�K���{�@@���ę ������j��C/��MH�� �0oi�{7Έ���{��)�%j1��T�;I}��1/���+��V��q�?B��w|��ַc��|�j�\^k�".�'��9�H{Uz������-�UOd~ލ]C�K#B�a��qK�~�I��y�����6�SSI�~P��;���Cp�6ކz��������g9`v�#�y��-�@��H�<)��v܌K��[oR����Ӏ`X�,�N�ƕ��5���pi�]�Sԑ�]���R&�F��B�&w=�5�&i��yMF]��{z�֭`@ ǚl��.�%H6),��*]F���TY]��ø7�o�Z�3�4�3�(.e�e�@|s>�5��;�<x,�n��%��?0&�ɟ (M/f���f��]吽�1Xz ���� Ou�l���p��N����hO0s^�d�����I]*}�5a��ѕ����`�,��/q�ǯ̿c8��v;j_Uhs���Y���j��Yt�#�G��������*��l��ȎX>l���+נ6|R�_$�W8�e���6p��[�m3��`@t��z�\��&��O�s�G=6�u���E7��@h.�#��tv����4ؑ�S
<m��V�R]�W��xd��uO�@���_�L����â{��V�ܡs+��EW?����m�P�_�^9:Xe����7jr���6-۽Cݚ��7ؕ�t�,t��i�A4a�2�|�����pt*˲���Ψ�
[wm/��������=�U���+w���c�l�ߌu��aQ@�\�'��-'k�U�MFf-�K^�j��i�T?	1�t�5�I�����Od�����]y��#' 6��Tfݧ����hISh��̝m��*�t�[*B�|�1����>/]�.����^�M�rO��ZqS��1W���� #��:���N+%O�)o V�n7��M�;K��n����nUzAj�`-��𐈙nT*M���W����xx|r033�G�	*�1'��3��ſ"����S��B�SH�f����|���a��9�r�2�;jX���\$�睎�Z���~��η�߫*W�*3�J�kmrP��ǪIOWE*�'����6��G�(9O٦�MM�I'Zz����l����,;i��%�� �@=V��^0��SZo���$�T%SԪ�#���W[S�ǌ]�,��B�>��o���EjP�+b���-��h�
��8NY6\�%8��� �9��̕FGL���<�2RAֵ�=6���e�?G��Dg{�?<��U�@��g<����Gt���Gs��'���5��wǣ�G����I֥Z��i��j]P�ɳ.�����w蛔iC]��U�Yo�PHL�Ǥ$R2�O���]�>E��p���@���L�{�o�*���z1�Dد�SǞ�Jn�AH�`X']2ha|�5����2��v�D��		�_F�#M �w��Qk��qa_8����k$��OzC�Uhq�*��E܈-��5�O�{C:�5�1Y�ު�饶�v�Ծ9Q���Z�4�Q�����A�;�K�"q�p��v�H��a,�ݱLŨD+��O7�%���	�y��FE�?g)f�>�������?iO��*��lF�r)������/V�����ǯ���M.��f���S����Z�2 �S��� y����)1��{ק����g��J�_��q�����`+^v�h�f�bu����VP�|U�F.��\|)%�PZfkC-��B��>��]&��=٧���Z-h�ʿw|�B	P�v��WF��x���c륩���9��/�	؉�wcC�JK~fʵ�91d�U��S���I��-"P�6��N������/��<8R�5�$f�n8e6d�ӗ��?�9oO�5�����YawxVG�NTr̡�
�Ť��0<=&�%gw=E��d��W���+�-�2ōޙA�䃶��n;���j�
ūnb��RZ:ީ�X� 厊5H޶v�!X�w6*u���R�*�Q~��!���[g����Y-�����g[�����-�6����!�!�w��Y�ݬt�%��e����D9������`�3��j*��k��ir���&�.׼�~ǫ}����k(������C���Wi�!a����B�K�.� �g�l(1��M��=�
���a���c߾��f�:7���=O}w�����(�t�����)�NW�{�e=���A�<��ѓY���wk���`5�@�8�!")Gr-�1�U_��s HV�*3�L�ND*��Dw��\�Z\ӵl"ׅF[�6�-��hr�_�&Q+�A~��7��5[pм���y��Ck�R��b�ԯN��Ӭ��7V�Κu�XeO�!�p��j0� c�(���Dqi���?�ٓ��ښ,2��Y�N�N��UMQ��	|�!p�fpV��ˢv��A-�Ⱃ���E���4��L�mK*�����g��
B+o����$�V"�OV��p�;�4M����=r�,�R��4��#����(��D+�K�"�/������q���>{؍�C���Bx����~u�S�i�v1��n�"�����Ƿ0L=0h�Gxo�.�cu:��]Vdd�@Mϑ0G�U�44�Uc5�2�0�e�l
'9.�+KAu��hI�K���[�ۆ/]�+#6��h�D=�'~_�"�
�Ƞ~`�ƫ��=�Z�H+sh���wܫ����?u��m���Þ������f��͖*Z0`�"��{·ß��%���e���ﴫ��v��#���x���ȶa��,�F��a`�像��_��1L��:t�M�k���J���K��Z�;�y��g2�u���'E �8���8޷p�g�$Eêm�J�L=� ;�;�^'�_ł�w�(rv�3����܌ǜ� �d$v��A4M��"v19Qg��	O�«�9\)O�Rt�wO8�^v������˅k�/��/���	y؈X�t�k�L���f�l���O�M'Z�t��{�'F�q�h�BkX�L7�7Cz�h<)�0���-��ŀf���T�����H�HB��  :�b%R��c��cIf!h�A�����x�x��_�=F��5`�w`+�6�}T��l�� �r8��c
��_��[��Q�ٰl���4��y��3�h�N*b7m��x"���u=q�z��*��<�%�*{�
� �Ċ�AR�bR�!�sqn���y��ѕ��ǋr) �ۈ,s֒?��*j��BeT���T��	�(q_n��eF	�;V��3l/q�J,A��`F%wj���1?~�ڄ@u��I3|&7i�	8Z;�edߧ޿ؓ5�$h%[�}j�K �Уpv�κ�V��� ���hw��\a�KR���
#S{ؕ�4����˗PW'ϴ�;�x����lw�J�P�s��F�]�z�],A����f�w�jT�cq�����?��1T4b^���fĸ%oj�庿u̢�~-�ڱ�<�������/�cz}2��(��d�221����~B�Z���*^����I��((�8��sh��*���L�]n�dj�,s�����}�p%z�T��b ��4�>^�Ot���+\�,�,�,F9�5rթ��V�� \ȠAZi0��3�1�%*�h2C��s��yI��
�2M��S�6Y
!T���e{(� ��#ߦ�7ߡ����E�t����Ͽ�b�R���g�5�=�-U>5���^fP��6�i����_a���V�Q��:�J@%3�s'(5V5s��G�@���`���4�� �!0t*�ҫ�o���1�`�oLM{��-���u�f��F2t��"�I�g�(�ԭT�'밋��v��M�6^�����}��3]eBDh��6 5�2�K�y-3[۠�Nz� #Ȳ�Ƙ	4��7�\`m'>A��p�yoHfi6r����pY�MY�A�¥�hH�+=S���x��]aY�:~[��{(���y�:|�˥��/�EA�u�Yl����4�j�up�	���������s���IA�@\��K�B�.S,��Q�L�BUd|���U��:��5����d��Z�4/�g֨�d3Q��Q�:��]шB���F�ʍ�'�B���h	/F}�j����]��S��x�L8=٩iSzǂ'�'�D�{ �\)����7e��鬬�3�7�#(5LZ�6h��&hI�� jV��#��lU[�0���~��1�J߆���ֵ��;Uy��xK~�+�Wc��QAq���(b�S��W@��<A*�{�Z�#�v�;��\'��V���Hk��-
�%8'�ݵ��j�qH�"n㈈S�)Wa˭�aQ��_���V���g�+�(7�z�G]ޒ>�����~�[B.����;Y��h)�59�mA�-�e�I]� `�d�[��V6�8U��WT����#.St�:ϸ�� r)m�F����0�W��<f���#�+޹�2q �̉�	�@��!��pn{�����g�O��9�T���&�J��}����X|ukZ!�Z�����®<����=�'�ɛT�G���3�:r��� �8h�e�����U�
�0)}`aM�>���	��6�P�.l���ʆ�����<�����De�(���lAm��OnQ:f3�2瀶���,�S��� 6���A0l�����s�Fc���߹��fUB��N�biJ�ފ�d�.�<���5`>��gHU�L�sh=���!��yMԡ9���?F��4���i��3�}!K�o}���q9��C�V��g(��s�>�`�����efN�>k�?��2F~g��7!�	��}������A���'Yaf$�tA��zs����H�����j��Vږ�8�[Bng�쀤��.u5�9I(=f���Hm���04x��E�����Ըn��F ���2?M /ݑZ��%��@=$��֩m���n*����).��"�K�.O%*J�D@�!�r{bu�2-���%���0�M��R�p1v��ӄ�Fa��%/��q|�ס�+�`����K�q�ԘI{�G��<�mCqHd� �u�����O��P����ӰJ7w��@�@X��"5B#[,�P'Zu�5�2�l��fWX&Rʮ���v*)���=9�~���kŝ�x��H�^I��$E藌(XV�_̤�B���  � �F���,ta��P�#e]�_���s�Q'[@N�5�ޱ����N���i��*��'QҦ�KT'x��ُ%`��fQ9FB����!FRwSC9�T�
�B!ݴ�.K%@ʾ{D�����aD��S
�%�Z�H�����7>Y�w��\;W��o?o�t,�d?�tF����S�������4�8���wm�φgR<�X{����=3?F�����F�ާ\����h��~�wu%���XpT<��2�`���겺u��`(4Ƕ����:AL튒 Z=����0ւW�"$�5Q|��47��m���3^XE����S��A�UL" �qj#�~���|�n�=)��z۞.��y��z+��#3� zqJxoh�Ij^/j5�ReO�g��+�kc�m��D.�av|r��H�?A����yv�L��k>\6��d�K{�1M����{�-����4��.e�$�W���""��9%d��u�3t��Ӓ�, ,��mV�7�#�����E#�ꦿ�<W�M<>
&f��F��=R0�Z��� ֌I�Ǆ�S��WuO��R�}s�`&LMi1�O��h���1U�������^�2�/�g.Pΐ(�h)�>��)��s4����m#���G�pk���x;���-��F��   	 �-W���'��d�>%��(�~���Vo��
�3S��0M��X5�g�t��`:>0}YB+��,DC�M�)���L�(�~İDy���Q��-)�2��U ��1qR�ldn�R��!j�1f�w�O���й�F+�i�&@ZI�aj���^��b�A}k`1@��^�bJ&zF@e(?��7U�?�]~r�r�<��}�4M[ٯ��y���u�A:? �a�eVS��L���C�x�,\��$"C���%1lh��*�����ֆ����;��~	�*��p��z�g�nr䃨�Üwm(�31,�b���B���)4�.evv�/��!¡�>��9�Q����7�4�y��c�H�r�&�o<J8N�nH�~�-#�Z>���|����&[�4p�����x*@�[2�h�����55��X��y=���7,�%�XT�X����v?��(�>je}��N��)�ֳ���S�Y0F����M�8�n)�ګq'V��1�,�%zd��a��K����+�hg��B�<��M�4OM�[�[�~�t�yj���3������Z�kG��9M����ى�Ѿw$s�k�˒Q���P�|Nk8�v�^�ߛYX��s.Ә�ݚ�+�U�5ujL���C`p=���w���̀�<f�c&jE��T�<�[���Ie��������3�i�v�����Wb��>��NȷP�J�"��{y��G+���j����m j�,ŀ+�C����	K
�{CִLB��wGq|��$Ƙ퍟0s�Â�t�Ӣ
'_�]����\� �"���PE���p�s�g�s��N`���nđ�nR�:�Ź�E�-�O8��y�������9(� �O\6ig>U��y���:�x��Y��8�\Y0�q��W����{�u�ӹ������t�
���T�bҟ���z�m�7"��qu���{Y_C����޾�t&wl��2>ҷ|�aۏ5Km�\��j�sk�r۫MO	�e�+�&�⪥�� =y�B-����9,b���Q�mu�V��i�ǃ���0ۼ1�)��|f����\����x9�c��ö�|&m\q�����<l!)��j׀��Kjso�D�9)*o]�gDOy0�Bj��yJ侮���r�
|�攋���ZhH���K<Dǂp��"�+ ��^��E4�>��U 'F�@}���ȣ��QO�����2Ca��C��a�M���n/"hrI ���i�?>$�:��69?1�3��NT�ؗ��NI׆��Qѭ/��w�%l�ke0�]R������wVu�<03`�Z��A���-@� �a�]�.Nu���7x�����G�ŗ�qw۞W��<ZVOB��	�tQ�Au
-�ּ?�;\r�,��Vǲ���|fR�Ѥ�/s�l�C�����x�N
X±3�TY�z_�a�@1s�6���V
��s
B+��(��I�<G��x*2���+��EoY+6WGbA�Ӈ�9(��ɳvE�/�`� _2Z�m�d�E+����������!�릇B�PbD �f(Px��
��N(�L��?��(J	5���ipL��ﱫ�+�Y�Sh��8
o�+'��U��/c䚪1Tj�T�O�%�T�/�+%�^����DE�칑�)� �m�H�w��4u��