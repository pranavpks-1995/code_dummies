c#���|<���r����bq��ZЯS��F�ˍ�T��p|^е[��-,�!�.� ���u��Ə1��nRB-߼#��E(���M�J�����H��+k�U��#���5�G$ÔfAn�3�e���k(A�DM�)���u��/U���L�]�H�۫{#��'S�:��n3�bmv��q�	��e�^�e��	iQ��,�����<Jp���j��o�B��uc��N�r�fP���l�#���;�fTA��Q��
��BCAN�D�D�;���3�CysaM�XC��y]�Z�獸� �&nM0�@�r�$���΋M`g�2�I�8t:���<S����썜LW�N��n�������dc�,�ȉQJ5_Yd�	����_�!��R��/��^�p�|��QH�rhiq�3$��|�zM���G|n�YgF9��+ �iuXB�� �[�_�ɢ��Ĵw��j�]���a�t�^l�l��%��к"�H�%t�����-��s����]��e ��{�J$�xR� �}+$��9����|��
�g@����	��D�|!�Wä��x�)�
�ό�mˋ0=�XD��Z�[�/��IEL_���	8��9�\�QC`T���� Kj_j^���l�?ZkC��yn���&[�<?�����M�� C�@ M��(�Ad�+��T�ޱ=@�>��c;��ʍh��9�J�,��]fl�s�����
����n�	�V�޲��.��uՠ��Kn9�eQ�oh�� �;v��,�X�?,{�a�-MU��/�^�ϚzB�)��6ߖQ`��]�Y��X|Ӑ��@~�2��A���P�J=���S�:�N��a�TJEz"�g���fa���#����@�NaiO��-20dj"=�-z(�A)Q����|���hʱ�Q̲�0;��M�ܬ9П�T%`�B�M��7Q���DD��L/.�0|H�{KL"�Q�L�:����g�B&��V����s���^? {Սk!�G��\�H����o�!�!3 �S3y�:�/"9����s�O��6B���^�m$}�4[d{��)K�̀�G�.ZH�P�}�BPW����@E�0�8�YY�6;}I?Dǿ�'O�Uce�@X�9�L�>��h��&�=��hD�W�c��_�*�n  ��+%�d�8���P���3��H6��!>g�NqU�)I����~��`�!�-`�}���LO�ɢ`�:܂-i�R;�t_դ�&^�a��#@N!f��r:u�
�~!�%��)�Z�J��%R�Yt����UٝcaK]�u�t8��;A�}����マ�'f@%�J��|!��:�����*$bNT�Q�-�TȻ�ٛ��:b�~Le��Q�k��8�]��.�q����#O�g�'(�E�2�Nv���,��1*a>����t�b�_v2O�	�b% ����U��t�����$M�k�T��ֻ�Q�=��'�0�	�k�Ҋ9��,�V��6��L��;�3cp.�+o���5.�Yp���h6mJ�m������ܶ��V�u,�>�Р2���^�h)i��./ق�v��C�Ɯ̿+`����5�b�1ӷ�`�{H &�� !�aL��e���ư�T/x|=a����F�@��R�1��A3�vmX,T%�OL��ےM���o��s�zɡ
�aF��6�V�T��}�[-B^���ϴ�&[ECᑮ�#�P�ag�&[ ��b�⤌@q~g�q��`�8�N�����2u!g���&���$�~{q�H�p��b"��ȗ���p��Daa�e�;}x����Y�8�Se�F|��Y� �{��(�X�1T�L/Pї���R�����Ѳԍ�@)���%�#�f�w����N�!/��^jm��ƍ
�p�L�IRpS���`���u%��6��<���^�Gd�*Y1��;WQ9xa9�n����a��������7�	#w�\F����k��g%�-ۨ��
jRP���}��F�#��ɽ��] ��z�ۯ�f�e�q>��\|��2Uv_4�@`��,,D�s�`��_�k8���8��٠������r�3[:0��k="B6~�逗����J����?�%�oĸq��ƑWQ�����ZF�q�=�=�H��⌮uh��tY�ˤw *nh>��Q�q��a]�s�l[.Q�܄'��O[G�{#�v���\��H��^>D��z�h�6���ᐇ��,܇[Z8���sU�`	�cW���� �����H�����I#�^;μM�e(U�� ��	�a<ڦ���@�y�5�l�!Sk�޿��?�:EP;2T�e_��TZ4����neq�����<����&�m����\P�pC���p�3Bo~��J��*ﮜ_H��~�ӓT��t�DD���33Azϝ`d��7ʭ}�(�ɨ>G_}��>M����lPb{���l*W=���B���b���3"���[�~|P�#ld����>�?(ړaU�!DbN��n&��kxz�����|MJ(�װh<��t�`�g4~ʔ4!��'Pc�\B��<��)����M6ksԤ�^G�䡜qa+*���TD37����S���A2�2k��^��>p���B�P�MSA����γ$cA`���/^�1D)��r�Sܨb1�Y����;�x~�r��k�-?��j��]�5P��������9hQ65>ނ06�g�8�Wѐ���#�I�v��@��̙f]��J�1B�K��̈́y�v�n����Ջ0����'jt3�bS@0�
Ik����8��K���"*m>�2`GX8��?�t�-p�.Ӂ�-��N�"��v��i�2N�5Iiy�P�jma��5�Q)��^P��=̐�c�X������C��&��=��������o��Q)D��A�R����3��X#�i�Ln�������!iy4Z�����&!׮;q<�*�Q�O���p73����	�'�殡��J��wD+�rM�}rb�<�p[��C7�.���-�̔��t~na��l�-�ͦ��.�S��ď�l=�Ќ'{�=��
 �`ŉ��D�p���	qh���X(�G/���k��#��aK�7q�sO�㴝;�
��Z�m2��Aq���=�D!M�@�����Ѓm�=���P-:.9�#�8�I6�$���N�m��$�J�`���P���?!�c�6O�xp�s̃e����5���0��\���p�`�ᐶ���.	�"B�ˡzU���S���Ɖ�]U|��<�-�U��#9���$��S$��Vh���#s�U�ym�B�w=��*��Y��4��ǻr�0<�߀���A �?Ym��`#�߃���P��,�	�����Y�ߘ4����u���'���2�9�O��F�t�f�3n>r��5��牎���~)���$a�V�U��@o�i��M"/��Ж�~�vx���X��λ���D��'���E�~�1�~�)<hur����ac[�t�(���;/jEYgK�o�tcL�a�O�C��m��������oI �}@�ϱ ]J!�}��0� �D�طӀ8n�KѬLp���Ś�E��=\���;S�*�;��(��%��:C%�w:���|�tZs��

Ĕ�s>�����i�RD��m���0S������Hq:�W�<�Z�Q���{�7f9�c��Z��R��¸�+wk���(J�`y�tGưT�����܍V���y�)F����:����u{��Rڪ�)��O��J��W���u49V_�n��SJ��	��Y��V,�ӤQ�L�J�?&�ё%���� ��PS��<g�͙��u#�ѩ��ׅ
RA��̎�Z�fig��i�4(Ğ�o�e%�����w�$�.�Qa}(,����C8��C���l�tXr9��,x�s7���OӐ
�ą2Z6�68ޚ��K����ڂ?x9Z��R���m������kU�:ɭe G�f{����e����2�e�>����c���et3�n;%L:M�_ͨD�e�t�9��H
�:�Ɖ�P��`��ܭY��lrl�=0$=k�{���0�`����� ��1��2����b�(�(QB!;�(��W�V=��_��U��W!Qih����JQ'h��2�ET����?���ƍ"o�&���A�,�c�,?� A�s+6�u��^��-�,�Ҷ��TCâ��rp�Z��L��,�W� G�,�KIe�=�������D�j. ��<�J��B V�᧶'��=2�A�݋�CU��EX�h	�V>��aƣ��,r��GH������^��LF��]OP�9��G���`�@	x�e9�k�j��jcYZ��D���ϜS�.���w�F��~ݭr\�J�EhhA_����N�pޕ��Sx�in����m�0�\��\Q$7�o�-2y��:��\r����7�w��ZGWg{��]�6�!�g�*M�c$�)#���+���#�]})ӷ��gH����de�c�B���
�o?+x�g��3�#D�#�{��O�{�u����7ψF�h�����/Hn�E��6��d�5�"�NFz�M�"-�T�P� �Դ��?<�NE�I�Qgc�sI6�n��/��Y���QE�V��ҹ�D�4O?�S��;�u�Ya9R�	�E&�Ҵ�s��X���� ,�S)�AQ���x�} "�S������5޸�����]��A+F�f}L��!��F,;����s�4#=�7�ۆ��M �^<P��T����n���i�n޾ϳ"t�m�jU׊�f�,��$3�V�k���8 O�����uQ������|�*$��7�@,��r�Ex�l��	����頬��,*����A/�t���YP���XEt�����mz�a��������	�Γ�T/�`�5����]��g`�d��=h��Z�(�$������u�-y�ƳT@!�ݳ��J�����s~�����J�zH�D:"^���M�4�ĒQQ�'�g��5Ny퇽 �j�|X��ޜ&�R�bm'M �/��@�J��8ƴ3�-����RyhG��\�V<e��,��-U�/���u�zt�U5	ܲ�:���ͯ-�TJn�-��=���B�Z��=�����=�tmʺ�ܞ�Xz/�Cl����0��n[����0`��f�2�0�#�G���B��ؘAV��!'��j��kj:�O����~�dj��d�������~���7���`�f=Egz�����Al����șp�;�2�̡^Ɠ�� 7���W��a�l+woD��+�5��8����T��	��%�(<�A�?'�R���)K3�)��?{R@