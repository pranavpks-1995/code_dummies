j�d���~%�1�@6qs�1���X�7�N�x�J�Y��8��Ȅp��-�U��܍5�S��6C_�@-�b�����P��O}��>�����kv�,�Z���X�_�-zl��	.��َ(/!
r[��B[�5yTON�w��e�*<v��Pf�#a����n�
�Jn��ԝ<*�SxZ����m���,�� Eށ��BS� ���>s^$m>���"	ˈ����&�iUg��ek�$i'd�) �X����4[&IfQk2,�R�# ]����o�Q1Q�cW�qC3qV�Qs˅�%�+/�A��D�lq`@bJeI �V� <z_���U�K� �B?Ҟ����-�k�������Q�Mv�I���6`�F\���oa��Ƶ�-�$(��2�f��?���r�Of�ǩWZ��]���M�7�.J�,�1V��,N��G����x���{���P/��r�}���"�
M�d��p��Ue$��Έ�����0�G �j̝��tL�
��tkr��֣_�� �Q �#R>���R�� �Ԡ_DWz1��b��0Y���΄���1��3��k��Wk	����H҃r���0*�Wؓ8�G�L�,��Y�gY���@�<����,Cz�E>v�+;`�SÉ�� ����Cr�q��v�8p\ց
 ����~[}qJ��B&����h΂�����o�i	��gԛ��bn��5��Y��|`4��0i`�C�g���W`�>�s��H�fDl�^������>ժHt��@[�N�tnta[� ���}¥�#J��Z3���̛��R������F�b�d�3֐lJ|>3�e�fqߜ�Q�N�T��N*�����Y�t�-g�B�]��Br�g�[ A���eX/}&>�Y���3�Y:\�ilm��W�	
��y9���!]a2�� �G��ݡV�8{X�$�l�f�5��-�`8���/(>I)r �Vp�H*��  " ��U�$�i&�Ki���wo�6P+�"��఼���[�Hb�x���b�A�o�_�a^d`�����ߗ�.b 
��#H�S`���lip��Cf�艦����}V��O	��?��!ĕ�C��%�j���D�]Kd�j����]�+ј2a�T��=�? �y&�+ޓ5ڼ�v����-It<�?I�qs�ě��Ј����0���PhG���;���KTz;&Mi*�\qf�r�9�1Mۂ�\Gv�$$�s�&w�w������s�	`� �Q�3�g.K�xghe�~;D7�O�R��6	�n���<����Jk�i�3xM�E��
�9��q��F�^�?��6_Y3���h�v���U�Q�X0�0_}��v�����	*ګ���w��1���=�/�l��&;�������e���zX�K3
���B��cI�~����z&o79>����[U�[ H61���=U<<�LAxR�w˥I{)�Y<���+�"A!���Ƣk:*�qe�Rko�ڪq�LzG�c��i)j�W�#���u�L��F%��d#/)�Ei�Sj�����Xg� u�+彼0%���{�P�I�-
$wYh��䴶a}���P�@�0,:���Ť�� ĄyIڏ�cb��bK���IX^>���g$�2,�A3*�!��0ҙ�I��Z�5����
7����95�B�s�6tb�js����W�0��b|`��Day��/>�w⊲�#l�~�����c_2SD��tQN����Dj]ZJ,�m��7���1��-�ʋ�o36t!�j�N���$];R�����;@�/R��,�B#]�;ϥ#꘍���0r�G��>�Z2]�HX�`oۭv�v?(@���>؈�y)�����f4���O M����8`�]ƺ���7C[x�<�۸Y�V��
�r�	b)Fi�X��D����J�A�fnʂn�Y��Lo��![ѷcH�'w_�A��c햏]�jo� �>���>��i��"�Q��2������d��G<Aw�$�����)����!a��%�DT��F�9�(ϡW��֧�JZB]���zB���N�� ��-vX	�	%@[�.�ܝ���*Ps�$v���nsH©zL�X��f��-�bNI�`/�"Ff,Ԥ`�Z��\�mvt�+�[�%�"�N�5s8U���-�Kշ���]HvD�Wm�Y�szW���K�K%�&x�D㝇�h�н�R��w�ʙ��CVK��0�LN�l�k]����pͯ㗊�