����?�Wˀ�ZC�g͒YȷP3Td��ֳ��|�Eq�P!��I�y�/	p���m0}ԯW�[���s#M?N$n�������+�k�u
�;RͶ0hJjD ޙ��DW(�/~����`�,��^������f��i�^[�R���w�ɨ�o�(�5[-��7{-�.;F#+|�F��f���k�-Y�gI~<�j�Yz����˄|��c/Lj���ȡ�a��bH~w2ԺC�1	�ڹ���uE��;�?'��*�{ű��{o7'Ba��b��ۜC�b<�����x(k7�@��� �H�ҕ|ps�gʞH��&����������%�,�ft�����h�F��:?�e&jɮ`LN�H�.=5�S���ԯe��>mN܂��$ ��A�6�	�y��e���å��ɡ ��T��a��:����6b��"�e�*��xqg���ĕ��(�@Vg��
wl�ˡ,��x]�}d;�ә��j8��]^�X~�$$��H6�u�vl�\-��Ǒ�s<cV�t��D���*<�a��*@�"�:�|��`Ǟ8G�-(��J��^�5�O�Yj�����7�x�,R� p,�uN�%�8�J�pM�M��{��|y�c�^ի*Ne
՛��ZO8����|�@�/���zxŗb4A�q�,��2-���^��!�gϩ$\�6�rMA%G����	�"2o�,���Ֆ����Ge��7�X[�s!3:rR��+ε�E�����w�X^H����(}��+��Q>��R�{��L����p��R�󒊖07�҆M�9Z��}}YS]�Y��Ӑ�I.���p�z�~b[�o
&�8�u�����\��3���f��ð��I�'B�n�@_�D����bʅ��2�e���쪄��(Q��̺B`Y��+���%2�.ܿ��� N̜�2��7�����~��G�ɢ:�'u�E5�G5@g)���3݆b��I߆ǧ�}ڛ���v2K����T�%�.�x@���7�I��U&��}4�e���u]���n�Pп:��2�T+o�+��p�&�@�CI�x   A ��-����/,4��adc6�QGiOz)[#��%���o�S�>űghG�ʛ�X�	dT���Ҟ*�{�s��#��]���xռB��
^錵�΅�T��Bٓ	x�>�\��r���+�v@������i�0�\���0��g�Z� ��BwĞ�O�N��. }���kn�o�lڂ�P�;M]���)�K��G%E4I$0��6o5��J��I���|OR�p��p����[*�}}��Bp�ꀅ�3��b��9�3P\�&��?�5�h��9^�0�oN��W��ʭ��Ii�HLĐ^�PW�����C����OY^����0k�f��ԹlUD3�����j����wW��:X�]Û���(�w�����ו4��-�Ɓ}��e��ů���V}`)?�c��$�f���$mj#��L6���H��\���m��^{ϖ�:ȹn��Y�v%���]�^{��(_T�{hm��RxE�9'!O �� wd$3�vU��}�.b/I����Z�$������ҙiء��2r��\���������v|6-a��J�Δ��N��C��	V� �[��k^_������[�|�e��	.&$ A��*&��-i��K#����G׍��J:������m�W�BG�ѨoX�.e�R�O5]߮ν.�wQ�,���b耯?��/#̓��>H�bͬ
��i�L��W����{2��mUl���өTOs8-`朲�ܧ�HG"���5����9�t*�t$���]��njҲbeLUp���u�t! �}�$�K[7�:�����G
)�����S�`�C�+T����I�%&���"�U��r   �֠����C����N�=wÏ␥8/T�~�[��8M����k��FL_&��y/�l�j��v]%,��&��5�c�]SP����|KFsB���+���x��x8bH����˔c(w���� ����k.p�D��-G�I�k�Mk�ܐb���{����^�k�6�NV��,ѱ8"#�H�7ݻ^cIy=8
�m��s<%��&�PlC �|�k�^�L�֑�X�>������Z�Pn�G���y1�T�������tmL1� ��	�O%{�T+{@���2x��Q�䍾C������*� 8k".��W�JV������j�
LO�`�e	����{�����-�ӯ-=͞u5���PRtX�7�PC�4ڣp )na�DE�p+S��b��f�kg�����v$do��'x�<	�;ߐ-&p5H �V�U0D�, ��y�-,hd�BӲ�<�mԒ���_e�X�+W3����s�=�+BA���Wg��9?�b���෩����X�B;c+ʱ}�����0ƜO��F#я��A>���8m�8=
sk�#��|X���9+槫C��3�y]E�f����[��������ǋ��l�10���哝.��q���������>��h�R�?�Y/�"����*��X�;��*UL�ŝ�!CcZb%�G�-{R����Xs���݇��$� �24b����ÿ���7n��\�\S�yP��Q�.�4[���䅖��1��L�x����2P�%]�n�}}O5N��������	���!o
�p ����p�\���Ae.�P,dӛ���wA��~�Bm���פa���)�v���$��5|��U�y�[��"Ţ),R�K�#����P�[t��=)(n,�'�q�����Q�2t�_�ߓ�z���%�������V��<˂nPT73M����S�������
+{dd�Ѭ�Vű"����,D*�7��+��̸��x�����k��R4�g9�[<��{�{�$�Dc�2/��bpFb-�6;V$C��^�DJ�s��&�.���#�EW?����	|�.��1h#��$B��v*��7dFu	��v�s���Ub�'G�;:K!,|�Y�b{���CMZ�f�2r�o�g;��4�o��Gm
��\��&�D�ӿ{J)M;�L��,ן���N	�e��y��@�_K&�ĳ4���0�c�t� ����s���?������5"i�|��Q�]�9��mx�w��Z%�
��|�������*Z/f�X iE�i�
c�Q"B�&�n��2H!rS�K?XDY�]��?���o�J��7����B8?�]2H��{z�94��>J�aE���N7t��*�k3W�ޏ��΃�W���h���*��43��Vҩ6;��e{)�L�WbQ���K�#��=[T�����鋆tw��du}TA�2j��9���tV�E�U|��������g���G���^u�#�)V"�;u��gv�'�И8��_�v-}Iwr��X�_ER��^��Wdn����H��.E���6H���6��/�TTV1޺%"���7P����c}�9x}�ԣh�p����j�����$�XP��Ӕ p/���t���<���,ݣS�,�!�-��V5�
�~^�7�P��]Z/�jLq&�(E�M�� �͑�����8{�����$"ka2���+JN��E�b�� ��#,�[mӗ��r�v��I�3���B�ipn�������R�$���~�؟��D���r�G�|�n�? .S�^���A5��w�e�im�~_�h�C�/TŁ��\�6�R���r������`��_�ϫ>���tV� ��G��X�I9W�=I!�ء���:��jīl����i�.}Q �����!��B��v`�8�{�V���ؠߓ������!�j�0)��g�@��Y�����U�����=��v/��TE�F�����ٔ����Ә���(�7�,��SȎ���/��]0 �Х�������Lu�ɦmoD3�A] �����0}0P�������Pc7�ɠ�9��@Z��|)� �a�`�Yc��ɰ+��8�P����@q��D<�2 ���XW��+�9��F��qnlY��������i��X�9��Q�%�Wqzm̓��ܺ���I��&��O�a[��B�E���F�$i�ٝh�Z��w5m�􊔰����[v�_�!���B [�����(�q�'�<��ȔJ���U_�y�uX�;K[Q�%��'�<�"�`�r�����;�9%�*����#�m����.!09��d�ؐ.%����Y��u��I;
r���^�X��n���3�ML�����7H��:��hV1>o�\Ec �$�b���V��g�p,]��+ҮFٰR}CިK�p{Pl0E����ө���vJ.'�=Ӧ�0�3 D+
X
@�P�/:�+}D��CZFo�M<2.Ņ�-�.3`!d`�\��f��3���ʒ�!�s���*nZ5R���Qp�w`8�h�������:u����g!�:�t?�������-.�a��ܵ�� ��s~5�:<rV��@vZ`=���_ܓ��&�r��ĘiݳD(%�<�хH�S�%���$bϰCh2�`��,F���k���&iωfD~��������h����IG9�\����U,��L�YSe�& <��p�(<)��0ݣ*.������' �ý�z�S�Kr@�� �W�E��ҠW�Zz��	@I����o��~�3O28�6{
j���+�WO��c�.�/���.jy�����JVݾ���gy��T�b�z\P0�>#?����d�v���Z�|���(�7�|����~��Χ�4���
Hߝ�A��:sC���cL'&�Ib��A���1"��[ϧ�M�H�%��'@�|���|��e�6KM�.�NîW_Z�-,%��?�T��j [��r�g 
�r���[~��CMG<dg�5�E�S�KX��|��^ԈȳE����Ҭ�5}��<�AQ�AN�S	��gڜozV��i{7j8r�� j�(M�����Gu�/M� [�v�-���u�0 .�!_�N�8?n�:dLQ�B!��@*]H�\���Ýn��BCT{����������C��^�_.��L��c�Zh��S���)����M�2���ކ\�Z�L<��L���"Qol���X��_\{�|���A%�b&9|�9�"��	S���E3����G�78��x�ͽXQM�4�>r8�W�QjR�&���rٶ�Lߒ*�^��U���ː���Y8ի���Km�xBd��xkhUZ��2z3;{���	F �96,U�;@����jd_$�CM�+��kwv-Y�Q[K�p\�mz.?g\H⸸^���O��v+���eйx�cw	b����-+>���R>̿W�M$��t�Tcޅm�\+�,�'������-��#7�KͬF$+,DC���6���B��'P��J���`.����{�SJ���y�����JƶG $P?B����z2�U�"7�T�JO�fu���#�$h��g�R���*�,�4�-z��5�\%�7�0����ͬԵ��A�@D|�<ި8 6V���eL��b�2��?!����ϰSz��5EWv��L�=��̛����چx��X5e�l��!��4��Ue��: �c�C���>�DH�o��Xf��;!ȿ����r��$m�GX=�U/�B���T2�P_�j�6�g�yŇʴ(5����3��qjD2�X�l��:�HFѝ1iE/�ڢ�`&�@E��"���09��N��Q�;�H$����r� ��y�<��:��hoWL�l^͹��;��wO���-��Yt{C��x��r���T{�1��q�4nS��W�|OC���ԁ (#��ބB�n-z��T�\h�+/]�q]jEY�y�-��RLS@8��ͺy�N�k1��E���!MZgN���N�C�$�]���
����g�X� �L�~��[�Iy�d�؈<�	��!�V�"@��i�x��r�l��3��0�n�eL�y͗�;��p�c��B��_b%mܬ7u%�o~�zd`'�O&��ཪ��L�F �=�X�e�	�«�k���-o���P��X�kBI�@��0�l27�*�}~~�c��oPXCIɵU��`^�d���L�;F�����i����Q��׆�5�%���Y��Ox��\��X��O�V�Ů ޣ���y�S$j���d#U^�.�E{�a���n�#(�#xKu@O^�����b�(���X��jM�		�����\��9kb� �A��B�4��t�	�xT����%8Ls�>�Ϛ�\]���MA�L��a�[��s�#�5ډC���!�(��d+�Y&�Ũ�ժ�j1v&q�%O�k���!m���?<�Xn51��SQØ���<,dt���;L���/G�	�9HE��`���dX�b�Z��mҟHGO���W(XPĂ{�N��g�Js*:�����	|!j��kC�4�?�E�F�@���>���S�7�!���c�7*Aҡr-��n/wv�==u2VjWv�����k�.(���u��3$�����ʎ3����Tu�}��x�XR7%��;��cߵE4����u��Qt؝*7�U��I��~�
j�b��U�F��P�#+;R�k�M'-�٣�q������HV?��v�k}��w�W��eL�8Q��	E݃ct��~"��KaA���gꅧb�6��n\�r�o���h,h��[e.��s�I�o�����ϧ��ٽBuA|�Z>��J�(
jQo,!�1�hx��J�:�T"�"Wv�}&�|).�V5�h�㖬_a�Z�A�I���s	���X�2gy{Y�ǔٯcJ+�1�BW��P C^�nP�YXxQ�[�&�˷;�*��Ҩ8��>��q�u��Qq�l�6s6��doAwֿ̲)������ӆ0��:"7��Wpġ�+�zOi�̓t����	fί��`/�~쀛�@���X��Jf�X��f�k� 
�P�u
u	co��k�'탘��������ה3�a1��=�Dx�v�&̳���<1�ׂ�]��u>&�R �T)���	=����a�F�)&�����K2u��`�Z�(L/Y��b�+���L��H%�Y0������=�~�U;,��I�B��MDZ���D�pGy,fu���m��N>3j��)���|Ό�抳�,��ߥ��VS���i���B�\�!aP� ����u���P�t����n��U�K�J��W����j��5��~����`��$Ӽ�YZ8Ϟ�ǆHW?�����u�^�{�������BX�(=�q|3:��}�攐�;o4ד����좪U؍��lm�0�FU�'���u���_2\�[��%�Rغ���<�x���|��I������`�D�  ��B'R��c���� /�G��:�XMD"�C];�7S6�:O$:���%��D�.+���>S��C!���F�ᆺ�G?-��˹�U��O����J���wJ�b��')���t��C�6wy��&W ��o+A�jt��A�D*�Ȱ�2&��Q+Y�bĩ��G����߶�򰅥Lj1@��Nbk��F�E]��-�t��'����*cl�qCHų�u����?��N�ޛ�(r�Ķ� �=�v��;�a��ӂzޠN>� �LO��W�K(�����,�ÎlL>��pڴx��x�ai�tV�Xrwڰҋ�!\�IJ�hej��Ɋ��A�.W�R���+�s�¾cN��V��IԹ$��]}����=�Jm:�k�	�x��������`d�7��bz��)!F���	u��/�i_杽�x�q�{��U���z�B��fd,�q��̗���(��A{�|�~�Ռ�!>�Jܛ�R���� ��;] Gm���_�썰S����ރC�(��GF�7��(��/�[~a�#�X����dUo��+�������ED�%�Ls�l]ܺ�&I_���Y
gM�'���*%D�4��й	�{�Ɍ�G�PI��"K?�ǒ�^b(j*\��tF�d�Uʛ��닫e��㼼J�S��XI[�L`m2��D�y�Їe����N�Ԟz�e)��l�|���i wV����]+ڇ���~����������`04胉���
v'�����DA����CE�WS7H�"���U��_c�jh���&��|,cZx��˃g���+�o ����hbh^�F���J�I�.F��ə�G�q�����h��_�p�7��CEW�K] ��VJ���{����1oY�B�tNw��a}v�
(4�~�X���V�$0���	G��=������bI�EipcT�m�e�1_��x�����cs�O���ڥJ=K��V�w�;ĖWQ��9
�2Kq7<��(F���(�{6ɨK.�KH^�����ɨ''d���h�A��I����$n���{T��8�L0F�-)�0mv�Q��Ղ��#�ۇŪg�1C�F�C��y=��S����ċs$���wa�z��nki�D,����>�\P���&�t5��D.�u[�X�CS�C���K���G��B��l3.X�����x�8�lҘ垲W$�`�6��xC��T��<D�2���)s��) �T�)H���2������/���D��   ��U�!�����H`���R�^���)��0qtj���G��FZ����_7 �Iu[8{����+��$Wq��s�ǰ`�*vʣ��N��S�ٺO+z��aN&��i;��P��VU�d�i冼
��NY�1����� �>��(��Q�aU*K)c�O�Fk�(����C��kČ�I\`�^�ζ��ց�SI�W�ea�s]�1ǚz��7�6��n}�Fm�,��~�K�X�p��~3%����7��A1�%��(EOwJr�	}�	�ׄ��Ȩ�E���Li	,e�g��QkS�t]�ڙyV�mXf0�Q���x�>vm�M����RT�9�y��>δ�����N ���+�d�	�����-@5E10��ل�sk��6 N2J�υ��Sv��`^4�s�k	�W��Bt���|�p�M�A���Y7�M�c���m�e^%��x�;e�ߧ�Ų���;X����"t)8��}h�ҚdP([m�k����I��bF�j�A��H@FQK;Cd�.tc�#�$�5��E��ԇ��x���y0D;3b*8�S�R��e��mD��Oa�����u����"|��\�{�^�V< {ʻir�@�!	e4�l}����Ț���&`��RQw�⚻u���S�6cء�w� �ً�zӊ�dV���м��w|/��u*�S��z����o)PT�J��c���^��̂߱���W��,b�Ip^K�0�#qgv�1��
��ڳ0 ��w5~Y��P.�� ?0��2���n(Z�E�*|�����Jw¬ J�Y��b��\t��������~�+5(���7����ꀮ�{���19o��7߳Q f��P����qFFue�#2P4.�^Q�g<�`��,�+r�:~[}#u]�,�P��=�R5ٯy�.4͂~�
��N���4�'1!�b��9W�d�?���P�l��X�p@h(�]G΁�9�ɜ�<�#%��J�j0�Ac5�g��,��a�����?�?}��d�����g��أC���   � �&�u�!QM�S!��p��n6����J��oO$�i�r�v^+U�bD�ۈ���cv0.���}�D
\�dU�`iw����|FaV,��4�-�uG��s��{W������c���.�TqW	U��Kڰ؎	hcûJ��Wqd�9&yFLP��(��:u(�<�@��ZŊ�ZY����yԹ3��\�h ���{ �;�q�f�S�a�E��������#��)�{���˩o��*G�=�U+��=zO�$^%lџ�]ɣ�Q$8��&��"��n���0����=��`���6��r�90�����o5CirFA��]A��z�P�!��mj�j-Z@,��g>=`��'B�<������H��w�tG1j ��������& 0��
����d��@A!\�
p�y��w@T�T�5,�c�4��=v'Bc�.<�<@����I��#�=�|���e!�9=��9gו��=��)�����L69�ʒy�!�WYҥ�R��N+hMC�?���v�c�H#��5i$�i����== �V����k1�%G���}]Z��s�8�}���K��l,�jx�m��3�E�᷎U+���-�.�b�-i�������:}�̰����7�:�x� ���c6d90��+c�.�QbnQ�\�dw�R�ڒ�a4�.���ڀP�iYS�?��e&��0� �i�bM"��G�2�曮��0|s֟<%1-�`3���|�ۭ��L#'8�Ɔ�Q�O[����c|�����W�ލ�a�g>]�^YI4Fў������F���x��Y$x��ސ�Ԉ���J`�93[k��������7��O�Y!��m ʄ��,��8B��Ӏj�7jgu���$s`c��oX ��Z�/2���n -�@wZ�U���.#ly����W\���5w2P c~[;$$��my�ON����B��H   � �b-����	�����E�pR��}6��3l�Q�L��m΍�G�D�R]}��  ei���� VB0B����S6��S�_��I+T'�s�+��]��a��c����^v*����c�
4� ;;�衄������WFg�Y�j\7
���sN}
$`c����|3�X8�R�}އx����(F���K;�7G�H�����[������t��{a�GZҌ�]�(<�x�A�������^r���_�O���P
fĄ�1W�( 6D-@��0?Zbz�w�����R�d.���B��+�;y1������d�`2���a���U?���M�k���rd�9��z��{Ⱥ6ߙܱm�� ��{ �V�]��˓񀔉��m9��C.�3��&�6$?��#�fԽ���dʎ��|�yZ>Mz�gab{��#���A((E�w���^Ӑ�)·B&����+q70w̘�0l�`��Ҡ���b�3�S4&��!�l���5���-B�~c&��8ӛ�B{96��(U��*�����48F�OȬ�L�I������o��J���0,�'�lV�ϻW�Ez8�hH ��{�xwv�o��M�G�x�X#O��5���.���2lۼ���
T��٥�`YP�������� sd!�Ȏ��ʞ��;�,$��֎@��!��c�1@i/=�ﵪ��;��Qu�_�����W��lDNf��@��T_f�o����S���Ν�ܸhc|�x��^���j�N.��E ����������!��0�0L��E���QQb�+;�8#��B����i��M���z��A��@��_��Q�Z���_�^Jj�g����۴�G,�P��|Gq���T�sL�D�Wk��	u�'�uQp��yF�������e �|�x������'yJ�� !�Զ��2�E㔤ƙp"A�){1�:/�d�/��_�� ���� ���@/0m��<�?����q���v��	��V�^�O��(������E���Ѡ�o��#q�P7@�K�`� ,�B�nk����!���f:|�q� 0�!���� l@��a(�@ f��I)cŵ3�����TJ(X*�)Jo�p������e�B��ؤύ�?}�m�2a_���)�ʳ���� YΟ<��@_GnA�ww��[�1![�C��f��	�_�C^���yc|�]��4��=e*��x   8!�ܶ�.�� -�  *J�K.�?#�:�����3� ���X3�#� jx��a���_Ť6%���Y���[�S�~	)��$�m=[�r~�Sk"����5Ta}]� ���`�� �� K��u��B��� V�"`D(��
�w�,�<�A� p!����+��#(��5�L�P���b�?$�s��p��oV�s�cr
�XHfkG�� �Qjq��	�.t��hDD:?��,S|k����cQ�/�çS:�+W�Lc-������O����
 2 ���Pݤ+ٺCs�s`  �!���"a!��*�e(�������Z8�C(чm����a?j	m�(*�H�y/c����*f]���ąLfM���u�l�T���)�F}���Ph�Sv���Fr]C�w�tٯ ~G����5�\7��4@K�C�����;�}ny�?�   8!��ȃ�#��c
(��h栄���v�Υ���)�j1�%y��δeb����w�D_D���S�/@((��@�f⒕U�F�	�*w;]n��D���]�:��	�%z'a�I���@ ���G��?�����+�_+гl�����A��t�u=ΐ�I���  8!���1TBTR�j��X�/�����r!�~V����C�ӕa���s�#���]զ��k�zH�֣'=����"�N���FCO^� �����`��9$�ö�4��NS�QPM�˯���pA���u� ������I�m�F�)�{�:_���ܮȀ    �T��   ~���U��D:0R�8���`��JB�,�엵�;�z+�XqB��!��Of�8&�\/�p�x��b�Vީ	GY�62��.���e�R����ɞ��"��C�l����Uu������IM��	�� 4��)��q�H������z�S��o��=�J�8-Ke���P ��++�m8��<��7*���ɪS���.-�&�2����GF*��J���6\(���o�QKcF�d�ܸ��l���0� �H��=NK���*,� "Ж�Z�xRu^Qj��]jŊ��2�D��#B�.��h;8<,��=fn��T��
�l����ߏw�+��! n�"�����t ��Jd/�,�d�!��OKKpP�7v��yn��6�v�X������C2�����t�9���_%�VhE�*�a���j����hPk���T(�ݛ>�\�������/����	$�L�NˢN=�Q��u#���ԏ�gv���9Պ�m�8W'4�AYu������ k�H��������@q���Uj���ߪ`${��Ջ�|UR����9�ʰ*�҂-T�c�}�x`�k�>FIz�w ��������/m!�fX2}U^��)���៝�s|�R���ȏ���GQ��Ki�~vB�=Ӧ�7s��H��������L0��ѫ�9��~ dr�_%�uJƻHt����O?��Q��N�Y�uV�/g����e��(���6AZ�K�َ�ðuF�_]��E�]�.�0�2��;��~�=��$�F�Ia� �h_�xw�eֻ����Ĉ�����3x�%��!�`Ces�u����)��0EP�s��6����n]i������.����� h&p�����08E*ڻT�:T��kB%������ѧM����[J�$.�.��X� U�l��ʗ����-F��p{���p� �b��=�-�u+�x����>=A�Y��y�\�'(��{�\�2-�[U�R��_�+u��e��n���*)��a���'�2��u��?��ɔGdu>bv��"���XP으�e�P��̶���`Z<����p�ϲ����$-�f�
v�r8�Эu�}�|j�Y���[n4�����"�ݞn!aH�_!��6�l�3��[꣍�l>p������< <
�^Y������ľ=���X���?_�
�_���L��t�q(��dw5�xJF�J{p��*�x�ё`��JUO�0]v��J�& �ʴ�:c���oN�-���t�{B���(�)���G��p6���E
�ӆ�>Z�n?��M�JT����j�R�s���R���H�]>[|L(v���"�Q�����5b�[k�;͸���%&N�2���ܻ��1c�q��RtӾ�����cDá?�X��W���j����J�5#~5_u{�qFi��2���3P
�\����3EO`ek>r���1���KZlŲ����,�����aBp��y؋�* ݍ�3j=����u
�t�����q�T(q53.�Se}�ޙB����J�J�Jr���Uz{Q�?��, ��f�t��EK���cwN�_a��CӜ���{������Xj�6>�ܻ�
z��E�O���.�<�1~w̿y@�����ʄAs�
V�L�tv0���o����-�;ı�'W!�Iܡ�C`їs һt��������46)��.�/��V���sj�w'/]�@�k�P<v��̓;�`�t���7�b��
����=�bY5���n��:�B���"� ft%	a�a��kM�r��Sd�����y�L�����9�YM`�Ņ���쁉��)k�Q�Y�>N%9�Ӡ>P�]���㘉���TۍK\^�4�j �W)|c�3����j�������i�c�]M��M��x��@��7�a� �_�A'�
�R�.����Ͽ_��v���g�����[55��Zմ�t�u�TI}v@Ԉ����@ �"1�)����.�{�����J��fa���9Tؘ�ߥ��p�!��B���xn�q�Y�0��N��a5D�vZ_ʶE���ngj}�/ω��Ytǣ!��[��_�H�Iy�����e�Xp"$��74(@�C(���۪Ym[B[{*-n���G#�z��6'����1Q��+�P��l��C�-�����!R1hk��_4>�#$��"��e4[TT��q�p�m��7/���/V��8�	�8�#���n�w��HWe@j/IN-�H�޺���صw���g{�����ht�I��t�E��ЃNϸ��|5\�G- �*\s��4�����i�ǿ* �l���F�\^�yV�@t�d���!��~*��m��ykg���bG�aN���]��G<��&VȶWwC���Rs�`��Vsε� /��b�aoD&��.H�����w���c	��]�co:�LR�����_Q��2�>�Ԙ��O�!�������������i�����с5s7/����Xj~:E?}TZ1�X=�Ԟ��&�E+UՏ��O��H��%��F�C�L^�HhmB	Vt s�g��dQ�xf��^$�G���eH��	4U2o�+-����x�����V���}"�������iӻ���g����:��n�����R6��Zaf�l@�6���q[�8���EѰ�G��&.�<z����zli@{K��(�b���2��[W��Z}ǽ��X�}�zS�]��5����)K���s|a/�'F���n����҉v~�9���?ۂ]�E�sJ\B�.L��N��sJ�C��pt�(���R���y����Y1g84H�<v����7zfoT��yAת�&�sP�%vՈ2�������?#���pY=� ��2��;�E���6Ccvw)QAA}��}g�f��4��?�V�q_��eH4i�u��߈[8�.��#��Õ����ʎ~���y�a_�����ӟ����P��j!+�6����7KQ�`�/��Hk'�Q�]���s�4��D��M��J���ʳ�*�9��Ru�.BAH899"!�v�!R����
M���{�.�kKg���������Ǎ,�~GF�v�A�L�0����� ����y���.��6_X���2a�>FE�b«�3�a#e��oQ�61�-��l�[�[����h�7b��x�Pp�TŽ��!�.G{�F_�'�&�����fOuW �~��í��3��YO9��ɾ���	��I �<�o0�"�(� !��%+r��n��"�T���:�=�}"g�,����ZNoJ^� zH��jn�&F(��1$�A�^i��V��3���IL!Ǩ0NXM��s�e�� �Q;^f��8Y��9��L�#���~�}t3�4����6�!q�N�a�(Y��Pc�5��&�q�)��\�������o�/f��x�G��,�P�؂	[7��F5{]�}�k�|�*�
G"��
;V/�`l,~i�|�wjV_���>�vĝ�+��B�e��3K��Q\�|�u�� ,��s�Mz�i^e�nOY��
��}�x�)�S�L�p�����b�iP3�x,7m��%|�x�R�"��JN� +p��& �@~m�@��d�#�M�oE�y��D��b�>h��Qy`Mfl��:�b�g��4��|�f��/�'�����9P!��S�;��*���3�	�s��c����Jw�
:tW�W��;>�-?�8b*3�k�75`�\b�ҪE���=�-�dm?�A�l�
�w�~��ŉ��F�VEx��?#�F�sG�)k�S��U�&�6�"~�3:�ɡ�5���/Sk�*Nt���1�\h����e�I =�K�����L��j���6Pΰ��c�� �1]�1���hR�#��$�j2Ť���'��yhN_9)R*sQ��J���]U3I� �MU�Z��:���Cl�~e&�X�l�%���$S��G+��85�B
�}9y��gK���� �~%����8o��T���HC��oz���z�Z!����<�Ε�N�`OK�>#Q��o`-~��^`��x��G(�j������vA�uG����ɻ�:S~6�{��_�H�5�AroCe���1�P؃�u_����@�܍��GRi����*�H�B�З�k`e���E��t�5�<��{Uُ1	�9�ݎǭ"�j�m�,�rP��͛^(��n���}��5_�Hh�6򫚕�X�]�#
�Vx��C�Z�s���Qe�v��F��$y�]��,�H�M*��V����vw��ڂ�Fv��+�[o4�S��Tz2�Vg�	���sb�퀴W���kI�7n������y^�������{U<@�~�@�(��3��ϔ6���nC!+<�r����w��G�!d*5�%��l�pz�`bC_ƃ����be-�����W)��4@�;W�T�����b�6�Pc��/�בk#q-e&T���?0��q�8���� Y �ˆvf�ž����]D#X��,ƥKg�C]�.���f:ϡQFq�_䮔{������{�of����酾��gA�~KSF����v�:y|t9��]����o��eu�W�@�����I�g�?v���8K��qµEΟ '�Jy��܊L;�ɠ�m�����TYG*m���8��ڒai�^�KD��ɖg�OtHM�Ύ���%�2��[CVW׍W��*T��d����#���@s�0]hC����6��%a�'Rrsd���n/OfEš��|9�<��oQ�T?P�k�sC��ɽ�Ico��D�8���2��oV�v��Z<F���y�)�mo��S6����H�k ��y�ꏅ��E<�f���$m3�	��ʃUKR|�g�Q� ��ю�(D��RD�Vx�_Qs��uAN��gR�����s,�-�k?o�Ah�i���Uk�����˔ں��Wح��+ݖ&�K���̈�5����R]�Gz9)�^�!V��)���A{u\�ܑ�?=��v8NN���8R�ݠ0�ꡄ�����E������ש70ɦUO���z���bi�u
3~�3�ab�bo\6�˂u�4%��~ʻB�(m(�����CqH��ϧY<|�d�=a2�
�9��^�g3 �� �5q)�=��
�֌�E^�p� ໭s�K["����amg�.�o���+��=���0eK㵂o���z@����d��'$�A��E��  ��%R��c��	k�ܑ+
G��:6��I*a'%p%0���Q����f}�P��~kV-g��l֘J�\�ྫŮ��ɣ*~���7����)#S梶��t��\s����'��&"��}�9�f�I���� �f�0o�� 4��-�1^�q�0���;%!�*�y�@	-"]�C��R@:��T]�V�>h��6J�|�A9ݿ���H	�H�5r*��RC��[�`h�kG�1B	�.;��[�+��H/����W�Os�C��G
��1��ɧ	�T�_��h4�'�I��.1��Tdc;�-�~Y��=L��i��Jv�!�R�QE�4��V����X�����l��� ��D~�s��F��ꀬ��j�-�'��ڤ���W�T�hE47�'A��y-@V��\�?H���r����k����r�Z���.���Q���q���aP9��l��e@d�����t�����'�H�R_\F]ϕ��yA��n:klګ���.h�"|���/|���wGھ;�������@&y֐{�ǩ�{�����(����b�oo�=�(�s�9��`�@�̢��?ћ��c�����v}l��bا������k��\6���� K����
��dv���b�*���oyzf�0B�̻��(9�5M���X�Aa_.$������4'���Oe��M\���.�md��O,�ڢ��zy0�Ň[�4@�
ȹ�	O���P����͆��)��P��h�@��Mh����s+�ĴC�_euD�`�Lk^����9���{�]�+��Ԁ����MzSX�DJW`��ɑw'��dw��Q=�F��AڠC�ܐ,��W��}]Z`�_+\]a]��~���e1}�s�/P�����gx�*��ޛ��E�,4
���='��%ݻ-�U�"�b��?� -��|���U"wd�γ�9K��7�@O [/\�$3��s��>{��4��VX�I�`߽8�w�?I��K	���� �-��G <.�`y�uO9x��]��!^�
�c߁1��k���͓��
�ߵ5��$̘J-���O�+Q���2��j�_w�4��S��͵?�u46\��ZWT�	Ź��^uh}B�^tv}͸�����u��QשiO^�J[��O�P�`���m���Y����J#�IJ�e���"��L�M��X��<�)���l{���BiKll�S�.�|W's)��TP�@SՃN�9`l��;���Wd������(^6s�h��V0
���u��y�C��N�[$2��B���  � �����,t`���ԁA���Q�
v`EH��{�'+�؀�jS4VZ�S�t2���ib�B�u��9�l�pj{���`�O�ȘW�2!�G�֪�-��f#�m ňs��x
���w+eʪ�,���Ť�L\�Le=��	;,ݳ�^����C�秄c�2]�U�,{�4<C��G����v�n����j�j*��(�5������،�_i����#��"�θ^lI����h��G�Ĵ�T(�x�� [X	�Uæ�xs�(�m6�٠����-Q��i�	0�*���/����68�H��v�� -�p�X��l�z��_�y����cO��p�gM!��)��r�&[��XrC|�[����^��&��u7�e��S��P^�o����54�v�Ok}2/Q*���t��B�o��#�1��@9������y�HP��<� ��/�d�hv��w�o�i΢jܢ0�D�칃3ƉI+nW~���Em%߶�e��ܧ���j��5�|���&fL���PP$A�������Noy� ��m'0*�UV08�Z�p�m`����}`��t#RM��B��E�,�����YC-5Қ�H9�Y�M��F|�0�ߜQ�����6�k:\S?�j�j�7M�+�A���   � ��-W��ã*y��冑4N6�Q@*����S!��:b\�=���!�u�y}�wm�M`�LRW�;���S�X��N��x8�bO�����\P#�;R�ߊs�f%Y���C�� �-��SٱƄ� ��n�3xq*�%>cBЂ�u��?��g�Fa��x�����[�B��!Y��%����,��~1��`X{�.)4��ַNQ	&��uӫ֤ �S�d��E�1��K���k��%b0����f��!H�Jda�}w�f'l�ߝ�E���{C��"�~��C�S������$U �r�}8Í��ߚs�0�祺���*��r�+B[<"S�!G�V?�w�-��U�sw���d���#wrGd�M��"(�Ш:�j1��m���</�먙T�Ě@7t04�XpoBc٫�r��r��]9�(G�.�)�[�|�V���   ����W�C����o%��X��䳬���w�7\Ef@ǀx�cF� @'�߹]��*�~��B��+?Q�:d?~�6U?osJn}qI��mMA�j�`s:���(���%��\<�N�u��.��jX�)����t1�[(L��8�Jj	�IJ`�I0�7�3��],��X�1����dk��#�V�q=�$�.io�� �K��|q��թmH.*��l˨����ۣ��^/�[$ې��Я��-��6����$V�CB��D�����R��F� )WYyI��&o%?��1f�z��-�*ZM����MJ��ײu��F,E1t�A��{�"��� ��-����0j�)s��2�}uO�gdw�$o(��x�G�$��+�c�&q܎�ո9@g
n(����y�����n�h!�����e��l�K�o�Y]�Na>���[������ ���TU�@���q���[p���F��U[6Kډ	����5aQ3��tM�:m(�7S%�S�'#@q����ܶ9�����-��XJ."$	�S
��~��&
�{�Y5H��%v̛b�=��=�%5�=�w� ��D �~�o:��@C]-4`|��B�J�<�2�ā��yR�
�͹��qJT�Z9�!��-oHʫ�hc�O1�Q���/���-f�2�+�`m#�|m�]��G}Yo�f�k����Ch�����n��=ZS➫t#���X*�W�4Q��->�/�)R��č�yV�wqHwjL�[���k����@W��Fm��cmxw�=m�������.�oC��@_�\���KH�����S4����.z.G�
����{'��P�n'����ي�~ � (�8?�v�p+ޣD4���A	��ޗ#�w�o���i~+��az���� �a�m򻻏��])>Cf��
���A|_2��("!���S���Êo�0��I�I��&N���3�fDRb�8�h{��bC�3��E=݅��c�-���b|��ޗ6N<�f�S��a?J	��C*�b&���U�Z�FzF��f��`��i�4�re�-����q_J� d�uk����o?R��>��%6���FS��#y�dj���~�[�o���poN�Ke{K'���^P��t��v"���[���Q�Y��t��K'�p����Y�:NxK�1G���W������?>O��^2��j-��zӞ�[s��=%����������Ӹ�r�2ݣr��!���t��e`��dM�zk�J�6o�9p\�ɻ��PՂ�f� ��v͗t�:gq�et�0�w����F�	4r��=�(rC����Ŵ��!�^Ҭ���CN	{�ٍbc.ѿ���"���q�8�W@�d��d��T��t	!�{9�`$��@�:�q`R�N36Oܗ�K*��iD�����7�:��C���POP�`�I��A$�E)y%U {s�'�N�q`��ک�!>���Q* �C�g#R#�v�Ml��|���F6mA��j�-���7���	!ikt��F�� �~RK��	f�+�.Z���\.�ɜ|��;Y�Η�����[���+����6�1�.=��>:�i�]��#l�v�7�L�MEYƒ%M%난��� W�@�\��Ɣ��b/�Q�8׉�ő�������o}M��7�Zcb�s6H��G D�[B� ��'��	O

�^�m8k�W*#DܒǪ��?2�-'zP��/���� �s�J:dR��y�d�&�4�6�/�1f.��=�ri����"�w�Q�c<j[V/r
38o���!�H����D'��Z;	�{ZK�5��t5x��������b.�;@,bb�p�֘�E���e���_�s�
`���.����0d_z�o�Ͷv�FyX�i��^pA ������!h2d�v�*�y]��!�%�.O2r���A=��oۍV�^���s�
�YD&<��5��O�N�\��J��JDLK�PK뇥���	0MKr�oL�IFqx� Tf����Md5( ���vSj9%ʈ��*4@)��0�lruߨ�m}�`\�i�>�)Y�Mbw�k##���̀ăPۤ��!��7��|í����o%{v�V�0?@�/�ç��t}�,,��sk�Z���6o��7۵�I�v;��d'�	�W�w& �<i7fBtd��Q�������r�AH�i����Ї��U�?v�����Ix�����JG]���ϲ��K��qĨ�YՐ�m�e)x^���y�SZ�Ok�c�d�GuT�c`!�0,K���8y���b3�y$ǁ	~�ӡ�'t�����RcL H�.��ճ�O�ɓr�+>�G�b��F�B.&=���8������qx��Bf�q) ]���.x����y'�^�0���֩�ο[�h.y����@���r�����ͱGm���͸�4�����U�
�@��L�C�F�n����А��Q >���F�6.=b�,ͭ��ޖ^��e�7��P�>����SI�����`�f�,V���+����dU�ߒ���;37e��H��cG�'1��w�� ���w�4!�U��a��)� ��*]}����_��2�0g�:�R�Ϡ� �[��]�`�ڌC��
h��zj��r��T���#�"�C���=�_�����,G#B���5���z#���0A<v�y�⤐�􆭾{�e����E�ezo
��h�7��A��wҞ�b����*i�(���cg�M�1���J�	h!z"�ێ�I7}�i��p{{����ϪH�����k���'����qxb��w�����V����\ ���İ{��umYa�ΐB���aN�~�(/t�8
�v'
ʢ�q	$,�jѽHצ���s�&��t���Ly���W����[F̨��}��"�Gf�(��z���`�QrB����=��?���������O�|�2zJ��"$����d��)�7y�
L��*Z<��l�D�}d(`��!��b$7��AS�ϞP�NqS���}�K4���c2/�H4F&D�f�G h�u�ǘ+ޜ�����)O� o�F�*_.�;�l���N	3��P��>��O�r����J��I+n�2ȋ��஄�
�V�����e	(��8��7a���!��D�z}a������||���#�b`�r����yj\�+xx�����H�����[����cE��Dɒ��I���T�y���/�wSNV�߶9���ݵ!��:g�j�����ՠ���!D��L���Ҧ��ǿ��~�9C&äH�7�:��H�/K�lR8�y9�yGv��}o�YU�Vd �����|k�]�|n��3;����Ë �[Ńk)tT��F(/0�{�\2.T(�L��J��;R=�_�:Z�]%iXA+T�v3���t-�(�l�QP(�J�2Ι�D���T�����(s&�(�=��\��ϨM�%�]i���Wmy�-,^_����D��t��*^�w@`#�$J_Q�v��!��`�h�+.�$����Sx���1���qT㞚�b�d苬�M��@K�R�D�E��x��'Ǆ�a]m�@�έ��ބ�@s��=�Rѧ�=W)��IL�M�|��Z�ԯ5ӹ�5g�STyۥv��	�
��܃�5�aW�Of��exT�ִ�r��p���N�W����b�&R�n�Dit�V��K�׈���#�#�daC^#��/����6̘8Ќ`��Pj@�H��X���uTj��ڌ�P ���#Y�(W~+I(D㒧&��ևT%}5v�Y��gV �,�������RZ
�p��2�+�*�n+���v�9=�TTX�(�]�9��P�FB���9`il#9?��A��?����Y��œAzC<a��6��H8���4���v�K!�_v7U��[Y[7ؽ����d�6�W773�zkY��A4����v�8�1�ȵ�Ǝ��g����X�s��[�@sq���[���v��o�&��U��q	v�s}6D�������Ŀƌ<+���Ia��P 7��n��-��:���t��4';cF�m�.ԋ�� �Ew���@�H�O���1N~I�2l��&P�I��t5,`��ى�ӮZAk��������>�,��W�X���8|[��T�i�u�ű��`H���y�u�ߜau�z/TT�4����9
���0�}��ALx��3r��@�t���;=�Do�(©������)��mDoHp�V0���Ÿ�^n\$:>�6�Teɿ�~�>�ꧡ=�o:w0�n��=-�Ty#��qs��Lo��<$+i�Q�0l�5aѰ� ����lW�>I�7_J�	S���H���d{�k�d��f/#Y�PDO�q͌���g��h�8b|�i�.��f�r�j���PqH�lL��s��/��f�ћE��*��M�(��ԀY����h����8ѫ��b����~8��	f�#9={3�j���7�|���o�+�pnH���6F6�H-�;�?�
	�2O��}v|H.����ǐB���j�?�1m�m<��o���(v�l�s�G����134����9Y�ӰAt�N�2�GN�_N����	��&O���T�z��N�)د�]jԖ��+�Ƽ�D��u��OkJ�׽,Qh���ky�N��ߩ/�/p�X�s!bP��H��]��_TT�-�Mk�+/.����8��M��TRj���;�>BC-!Ƒ��U@D�]�T�c�ر_��B���W�	�{�i�ۓf�ΐp��(]X� @�4�{��B�1]#|�e����E�ۓ�]���e���y�1t8��p�����jثB]g0
os��ndms�	ؘZ���q�6M����{tY��EE��֧Ҏ$�bN0�1}x27���^�@�n�U�I�aed+o�֙���<������۫����G[�#>9�T*{d�Y�w}N6rG��L�
�+�d�L�a��D��gn�1E��1��=��5�Z`���V8�**� ��2�䞠vM�KZc�x�{f��2���;��ۼ�b�G�@bA�n�����#�-4�FkH�~����c�����EJ��;y��o�k=֫�A_����Jn��L�k����h*U%.�pk�n���H��4Ee�Vɯ�t[�B�#s�L�yw���z;��:	˩|,��ٙn�[<��{����a)�ؔ��l�0�G./�����,;E8���Ѕ�y(=6c��¨��O��1���էo�����/;V��3#�IY�tR��FN*��%?^�[4e��Zp����]�`^ގ��亊��y �3!�����:wqp(��J���.	WO�	����"Oܣ���/W9�Y�t3Q� �5��~�p��es_W�����1-��"y���g�d����Z5'܊��~FN�PIE�DzA�!M�A�d"	B���uHr���N~�=���<r��
�;T*��C�a۳�<��k�L�Am���9B#0�=
��fmE�I�U+� W͙��/_��Fk�lF��g����Q���*��;cH�	.z�*��G�#[��țp���ި�?�]������J|�H}z�s�{ǂ�����Kt��؈`@pH���u��r��S���Y�n��[m�ǻԯR�o?����,� 4Ĩ�^}Q��2v6~$]�%��.o�Vy�/��#k4�9%��ش.8���L�kUq �viT	����@T\K�~�bm���s��LKg��l�f&�a���t)"p��^�J���-�Tf��6�3�Ѣ�z�e�&JRb�~�!1��C���  ��b'RW�c�#�-�R-��������.�3t�Mf���~ԥ�����M�!����.Eƒ��R���X�u��_B�9v��h���,��~_��E�����*���`w&�ҾO��L����%��ėn���j��o�>��jJ��p0�wM����1��ݠ��
�3_�]��N�K1��tW��)?9�}U*���5us��81���:��c�F�G{�	mC@��╘nTK�[ )9�AoVʂ:Ul�
T��,k�8Ⱦ��&kN|��D%Va<�JG���u7�@�����Zd�W�C-d�d�M�k�*����lPx9������l>V���_�bE(�2j�o"^��O;cO�R�&B�l����A�b5_����/���}@�sW�� x���������l��CWѸK�7:;&#��I���Θ��'��&�"�0���?��]`�-�s)�I�=.�^�a��S��Ez'��������� �/`=Ld+��I����5x
�c�{:�i��_&eQ-��=IK ����H�\m,p!�	���������k�lV��R�r~%�	����;�[h�r���^��{��t��"a@(Z��d���k����@�a;sI�Lbմ��}�f(_(�e�c��5��u$��<���	 �o]�;�_�&�tv[�65|e�qa�~�z�D��(E3��V�h�kw��in�U͝5֓��n��d�|H-y�Y�"yg�9E�˒y�Զ	�"nݝON1��'���dew��S��R~]�[�r׾ ��ڶ��a!���D*���!��@�J�q�<-P�R�?rhl�iǧ8 ��W�y���@��Y;Vx�c~�X�����P��	Y?q���6l|��+� �P��j�(]�Nă�m�!��_���X쀣B��B  � �&�U�|O����(��$}`�}m���cspd@��aO���2 O���$-��N����|75��$�������Čj�:�>����0��bE�Q��(�Ŗx<�Gq
���)r㈀��`b(Y�'�3d�OI��[):�5�eUdv�šJhs���e���7V��o�aC����D�jno�@�����U+a�%�֓�@Ү��Fl$�-> q eM���/	�<n+PͼD �L��w�L�Y�%��4�ދ?C�%�.H�T	=
�ք-�@h+D�k��x�A�@��f\ܭ��Fq�Z)E���`'z�{�w����8r�
���GN��T�NaD��g�
��۽�V�	c���]i��TҖP���4� �ܷ;�}�4���Ǿ��L#����ՌZ⚡֦Z�W�q�pܹ�ʂ�B��H���*�C��0��tٷ&��|��2�e;K�Dv�3�0BBR|��`���R���O����{ʣ��_���_��75/Ca�ޮȨ�4d�K������p�2��h��ȼ�?Kť��TE^�9Z��R4��K�����P�
�	�>tA�_q��{�B�_>���5���i���P��t����j�2��s8}��mX�3�8tg���LL9�A��S����ҽZ�BЁl   � �F�u�!\�u(|hX�~$}^=t�Y�d�M3�o�](��fYy�@�b���Hr��K�8*�?u��c�Ji�9�)A}oK�}l_K"�f��b�|���Jɸ)`Z1Z��Ԯ�P��t�ª�T7���k���?�{koJ�>
ri�\Ȋ��J�}�Z��F@�R�Kd Mz��F��[�{���yzl<�wn��{��G}O�Vm��kFP�	�%��w<������k�,�C�,"#�J�WeI�v�ZА��|�V,�F�Է�9y�H�=o��Ԏ��J�AJ��i̶�ȳ�E����5v}54L�V�zc�FԱ
�{gr�j|=hƄ~�c�׳���!y�k\Nî�v�"d�br��nH5`���xv�LhP����ԕ-}jt(غo�^e:��[,��A@A
f�}�bQ}d��dΠgd9����m)��%�B������O_00Z�,e;�s%܄�g����Z�j�1dFi��JP�Z�Ax#���w��i ?��QV7�pR@ߝR��
�|�H�X�ۆ/$�R5[�xaE�(���)Zu�^�9Q/�d=`����d<�^uk�!!v����K�N�P��1=����K���o63l�ojǲ| 
lq��Fe��b������]���8h�7oX<�O@#���eB��j?�B��.B3�h�Ѓp���ؤ���_���cB�|�Tn�BU��   M ��-�����y6�V���:R����XP��tY�V�#��E�F���x���Fq��J+��$��ZI�_��N�_R9<���z9g����$��|e�[xP>iO\��m�/rե��0
%���$���z�I�%��>y�?1ʾ��e�E���Ðce1��R�q������{u���L��T�|~􂕋� �U�;�0�J�Wb`�ZL?��މm  KVH�ت������"��@}@FD"�~gb�$����-�utl����r���\v���R�j1��S�R_�7$�� �����?~�^Sa)��.���>TZ|fD�ђ���ÿrֳ�R���!X]$)6��贩di�UM�辶ӷ�{����	�CF�#L��u�L����\mtQ�s��eDX	p�� �nv�w��P���r�$P���_�G��w/Di��9P��Z:��(����A��Kt�=wO�ʛ�����|��[��k_V�y@�����2��QĄ�btt4��<�ế��n��Q}%�-ׇ����C>�Y�@�`6����;guO��Uǒ%XR�@���1]�4m�_��=�`�E��	������ý!��ǃ���B�ڳR���Q%����"u�P4��u���mmKk��hpfД9Ђl ��4��8J�]Q-���Zu���J�ң�1Zt�V�aT*�ϸ2��X�*���L�3��7{Yv܅C�d�X��)�	�k�7����*j[�|Wx.���s�W:�:��p�0    !��%�F��&!�0���/V`Đey��[�Ǻ�����H���f;禼���5�ԕ?��ľ��U-\p|1s��c�X*�P��rh�?�g��hm��!εx٢/�������s[!����5����2�sE���o+���u@(B �	
3 FXM�"wZ��?R����A�$��m� �8!��=,aMՄX� W	�/����[�w��q�ߴ�% �����l�w)yP(|��[��)�?����@�:��m�M-q<��q�ͺ�^��/b���y���ș�F,�3M���Y�+U�="�WW^\^�<��蝍����b���
 ���|��^^_���������N�'�cnia5D�X%�x.���N�Q�H�@    !��9J0�]]Y�
� X M����[bx��&l�Y�4�R(���Up9��ӽ���庻�̈׻Ϗ���}8���ɝ�!G�s�|�v0T`���z�L�8fWO��i�K��������f	@���6U�`X�k�Xݱp����E-����ؤ�@@ �{��I�bD�]�7i*Uh�T��M�0 p!��8��$@P,  d!����2#:��%� }��ֳ�uk8�'LY15�h��W0�cOۘ�b���v���l��@*;�ҟ��t�P��ʦ��$"H���#�A�a��P�,H��� � )�_FH����d�%:D��R4\�@\�o&z#j���$�; ݤ*�[֦U���K@�!��=GCPe�.��ኄ���uG=n��\�7˕�l��yj��riQ,�!����KЧ�va�`�\s^�A��k��E�.���qF{�G�F- ����e�q�n3��-�hQ�9I����hw9\!X���b��Ɓa��pEY��6=��j�ŨV1$o��Ⱥ$�@¢����(]�%)\ @!��1(E�� K˭*�(	��Г<yteUh2�d�e:�S��B1�f�r�N�`YH2A��|�z�@��.�h>\`�j	K灧��=���d�p���Ih�KԨ꼆�������u��$�8H a X h$v0m�l�(v�k�����o��H�\�i�
����F*�AG$XT��0� !��8^���um cOE�d�O�Sn@���[�,������ۧ*���O�ӯ�c3&8�C)3X.���T
�`$R��
�l��p�N��~�i��F@B (aJ�@,W������%0B�e���5P��۠�XSy_1�e����!�)����URe֊����o�"6RV� p�Q`��   X�����C���,<�L��Rr�������G��w���U/s���əZ�OB������#�unw�U�~�Lۨ��M�V��"���NƄ�&7]$���a{�����d>�����T ����z�Ze`���fM�;�|�&�F�M����&�Z�����$m0�S�^�i�c�W����~���)�C��8�1]�~]�\2r�F���\��^mfp�0j�`e����h���������}M��g�����m�����-sᅱ<�˓w^�6!{�J%P��>�"n����\��^���5D�3��-Wpd[�\Q*���ž�$�dh�����sφ�Ao\��+7�ă}K������Zv5&��Tz�7x�7�Et�Ps�I�-�E^�x�� `������%�n� P�#W�2e��ɧ�#���M�P9kGY�h0I���݆NQu��ں#v񧩐m^�v�d�j;����"9��a ����`_�����@�A��6�F��>"���V�8qq.� ��F� ��\1��6{�6�E��	�>� !���#0\���-'y!_i�eE�E�� m�k�}kgH�x$}p#$��$uLs�F�����d�8����b��~��(�7tC��)�,�68�����\��6hI4�g�٩Ć,�!!w�Zm�l=�H����F����-U�2F��[�Rt��2�9b ��dՍ��6fo��yV���ť������>�]e��Ma��L	S�w�8�����E��wK����ϝ�u�>����`	�Ly+��w�ĥ�S�_ט�I]O�}FH ��(I5x}σ�¦�*�%zBp7$��en�&����#�����18B�<GrU3FS�	��9�5��=9�z|1�O��2��қ��&*ہ�4�pn�Ō�yb�b�sID��ݯ
���OH�\T��RC�������ig�uy��)Ml{ps�#U@��#ǫS%�� �&P0f�u�P�<�����:PN�i�X�dU�7��1��#+�ߗ�����o+/��N��0Z�s�`�fg@��e�^eìM⭇	K��Ś-ˈa�ȴA�������]&���b� Qr���U��Ixmq�m�4{`��X�e� v�Ějs���0�D�E9S���G�}��H�\⟽χ����ʡ��l�ˎ��(hW@&���%;x��t"׷��ɋU!�-��T�ϛ�:�v�aIo����2�����89P@�x��!�q�n�	�w�
+��;�	�IV�Ֆ�n�)�AN�+�YJF�h�e[bw�=�j�>�N_�e�fz�?�`�+��35[���0P�t� '�X�-�@��lPcXyx�H-�Qo$� ��1`���
�|'t�)��YF���`�M[@�I��)b_KM���{��1E��C%x�Ad�������Zv:g<��-t3��10z�!Z� �+�zY]�Vs=қ��'M���)q�����L�wAl2/R	��Q�;�ƁP}��y������a��.�{&E�=�ڴJƺrUļ?��- nҩ�)!	9��J#�UZP ����3g�?N��>�����O?{�V��p
B`� �S��2�^K�X��9�emÆ���~���a��Zct� :�@[* ^��m��P�#ݚ?^��8�[�r8�Hg��5vc���9d梌��-��ͪ�'��g
�ò���-ʩ�T��ŵئ��c�k�^�%��抓���+3�f�E�3Q��)&��I�"��McQ�`fV��S�4�]quL[�$�����>�ۗ���8�c91I�F��<uYGޡbۆ6�������|u��gd����qg����O��н	qI6�5f�>}c|m�{-Q!���tx���!%Z�.̼����DA��`nM5��+P�%�kx�kb���)��~�"`V�lU[��CPc�w��r�ŗ�������������G������)4R��d�ZH��d�0�h,5�JXV��c�p-�_�5i�	�&�>��6܋�"�b���hǿaB����:�aJq�s�v@�Y!���mM����$�L���/%��E�v�4���k-(Z�����'8�<�J)�ɯ(��]��[��JwÁx�t�{����?��8���C�=���^��>m\�k�9o�`�=���#4����A�T�	���������af�O�soJږ���͊��vפta�qx�����8ޫW�K��1g`OvL�؇ǰt�1;�Q�)6�d�-�VX��%U�.ޜ�qP)�>:�BE��P}���b�^�� ��`Q� Ei�~Д9��!T��	 7�`y9��i��8�\U�7��y�vʁ����I{��צ`∕1f4�|q�����{=t]�A/��[ڌ�~ӻ@��O�b-4��-��pC���T;�!m�	h!����pb��0j}�ݟE�٘?w��!̗�1�&(������}���#�7f�9�a9�Ƒ��_�>xq����gK�W���m�X>�u�̰�v?$�!�Ø�F3$6Y��2�s�ZP�I��t��:zz�|V\-�U{<<�8ɯa�w��r�$ rQ�}���Wt��艚 �T�M�ʱ���r�$��k[�1�)"��c�&�UR��'�ڗ�&��x�L�R����Ms~���ʾ�4����`m9��pŮ���oJ�$7�"Cس�����}�{�`��3��eg��Ť�:��{X�zK'|�%��*G��Ӝ=Q�s%�`_�PV���0��S��j�O&�ނ���O�dESM�b@�<���~]�� ȋI���	L;g��Z#?�z�D�{�-�����Y˜]���0+<�
 3��C@�;aU�9�h{�������	9+����r��̩%���@V��4WX#���mq��{���	����~��H���Y�Vr�H
���������w��N �g%�<�BiĽ���#���XP�Lvڝ�xQ|��2���-P.0Q�7n��_L�~S�v��مy�ʬ&�xs+ɫ;��T���V��+խMU
�ڮ��-�@´p��Ju�Bu�f�T�ʭ>����ȗn����@�e;�p������o.�N ;���dP�k;�;3�{�����Y��!~��='�U>�`��|Y&�T7��� V��bTF�̝�����h\�̖�Xgc,�#vC痀�˶Qc̫��I ��:*����:6
s֢�[���Ó^�
��>X5����k)�jpD��Ё��ݚ|-��/��EC�iat&�"rX1>���N��?���Wy4W�;9 qϾawB�f9i�.z$$��k�O��wԓ��C �ʥ~M��/����Xd�Yjs7t��˻����$��5��h��$쵗��@+g	��S;h�X��� jy3R�mrD�[�&;��J��`�� ��jeD�&D�|2���$:Qk���A�=��J"CO��GEs�v��".HF�$�������#�h��#�#LJ:�c�\��EU���# �C�S�r��D)�{&��R��;G�<l��vW��5���R��t&�"�n��	��v{�%�H�cs�m6茒fH���b�ml�2�=c�����
>��%��3l���𲏦��e�ɤ �I�tAݽX��g��Bm���ca�ƪ��Xw��\wF��fp�T��V�%��MM�n�W�8�@&�򜆧�4�+d�ETJ�����ևl���N}Utv+�j����gA�Fw'1����)>4"L�@�fW�&������ ٯ�D6�������F�x�W�<k��&򩔼�_��+AC���gI�#^yX8;�ly�����6w3:2. �P�oާF�Z��������+�Ǌ?:Gf=Zh�<Z�!�Ӄ�/��5�