(!�2IϨXj�W �9��m1�z�\�J����53��bd�>�,'�m��b���@�T�\�%�m�,��`��TăW����5"\^�(�=R
(��_ğ��:�N���˝��)���FR�ӍzZ�8D2X�5ƅC&���&�Y��b�uʻ4 y�e�*? �:c��5���9� ө3r9���>m��$���zԋ��J�����7�:P��潼 +�?�vk'cx�5ߡ�����.6f�����
z`r�R�z)��P���	ı�L1���B�Z�=}$����WaX�O�3gW�M�f����a?g�N7;)W��?Y:/��$���ꮼ������<Ԇ-a~��F������y��%I�e�/��Φ�ز.�"	�H�0��j�ԅ�Y��cԽ�֘ou��pBx:�\&`��]�z�efdfh�Q11���1ә�
d8?�r	ZN�q� i�*#�i�t7�=(��}�ڎL��P����0l�)����8����F�Yee�����s���g��3� ojC�/��Ҍ�A.������Z	���\bN�/���r)<9!7�>EB��}q�dF;��׼�+��s��b?\R�ۆ��`/Hp�j����4Z���� ��/l�6 p�l���[.W@�w$8�l�9����f{a��;�wy͟03蒉�QN=���1�����G�M�3�����|`�80��h?�4�-s�g}����0:0��l��(�f�-۲�@������K_?eKC��v�