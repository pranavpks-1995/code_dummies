Q�������a����������bq�0\��>  ����2�2s���_{9]�r�-$0     !��&Ca"D�&��� �/�.�x
b�-D,��[�o��ͫF3wy8\�5o����3V��h,��.�_���jԷ�o�l��2��*�\Z�q�E����9��5��j�Ls��6�,Yu�
@��F�V�l�h��	30| ���)�o�5y���Z�n��      �!��D��0�SvE���(�&P"ЬC3KW��%���k� PZ\kz�lP�80����q��b_��.� 2F�R��n�l:���M^�K=���D
���	�O �+�os�_ȩg�!�s�]^��{; �� =�?#����7KrI=�Ur�t�y�]��U8sl�     !��)%DD]o�ѥ �(ܪk
Aˀ<������UdI+y���.k�tO�����+�b�. ��%�L":֊��_]q��$5�n[�qj�V�W��;|Hw�?7���R��k?��~Ѻ�E�<��0GC
k
Aˀ<�����e���z9$���=cWɏm�f.��      !��&�"��XP�e��[�۷�#��KnX����G"'A@�=��|0A������,����r	`x�}~�cڈ�����O�*:;}�� ����������w
|�$Y�a�a�8�v���x� 	t8| �~Q���i��T����=���� `    !����� &�	�W�����(��y��z��
�B��E� �L�|Ǧ-kV^YAavT�H����+On�wo��`�� ���3u��t���	�SqPK������� �,�&:���m��/U��d %���T�V?�FO�z巃i���|�7%ﳯ���    p!��)�aU�e+3�4�,��m�y���%u �%��B �W�#Zf�X� 
�e?��c��.��{�  �� �� (�Ɏ���RĻwE�耐b��eYPb��[�o��^�2 dˢ��,� �º(%c6�m#7B;�Ib��۫�0    �MV�   Nր����C�����D�&�{��L��,��=�*VR-\��h��0��f�C�d\�F�{�qq�}d���La�<5����H�?��%�7 ���q��8)Un�N���Y�P��d@L�U�h`�`���;s$���Cm���9qh����0�I��6���	��\�m�ɮ9��3�?v��֤Tm��!���R�q����t+Is��bS�4!�P��_����R��U�
}p1٨�ܳ�*/��5]�h�F���o�`����61��wH���R��P�4�BUnw��������/���~R5fp'���(��^���T'�U�q���;�
&&�wwW�_��󋟹���˫z���{,)RPB*�7S�ֈ#�)h�x����CB�ݡv�~{[��Mwc�mfp�����t��pƎ��v�w�����TL�L��e��h��M�bH4R�K�!�O� 3k�!������[�-������?�oDm/�տ�������,hz�s�8j�,L36��
i�W���;V?�L���V��8B꤄���
z�t�4VT�s�<�du>q�L8��e/�̈́����d��>�ŉu��oy���fe;�[��R�K����%��yv^�ڣ�;Bz��G�;�zެ�W�l����
��ۤ�v���� =J����;�7�*-�P�K4i��'D���������B�b��(H�k�58�+	݇�N/I&bB)ԣrk�j�fU����~P��XҰߣ��}�Tә���U@��&����S��"�B��K��eΩd"�z�j�s�9&�X��'��h�e$�_�8��hi�}b�7J����Pq���E�뢓n �����M���{��`! �a1/(5�ES���!��X�m-�S9�$������g;ê��0>7E��La��ԭ�.��h��:��v����R(%�� ^�[t ����gT��Ҹ�ꨌ�β�^�N�/ܳ2iD�:�Xbp��Y�r�x� g�>Q��R��$!�s��Yc��c��uE�V�CI�k��䓉xc�]%�e�Kvs�(��/J����0�2�N<��c��a����7�aG\�Yx����