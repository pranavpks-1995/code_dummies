�Ca���ٙ�;;|�B������.�ɇ�6��Z�����F�`�*'T׿�}��:Z ���{��Hm��/��!恰���DZ��Ħ?�"�&�����͔I�k���ѣ����Ρ��Q�[�jم�l^�6ݓ���5�\P����1R5Z�UTG@_�T���o.�Q�	���ĳTw̆&�;_�W����Q�����p���'�ț�|k-��	o*���Yh~�����Ҵ��=���d(����e�B.�]y�E��t��Lx�Mh:D(d�ְCS�^�
`�"����f�ƀ�Gˁ }  ���xc��[/�VMDi(�EX�CN*v�R�5X�6��L�j%�`�i6F�wO�2.l�%�o��A��_�<@ԣ��Qn�y�seޓq^�eF��3�sB����9P��\�O��lcڒ�f�*�į�݋���8��HeC��V`�N:�`����z�M��v�O���tH���`K�}�c���w���6�g�Yd��s�<h�H���y�o��@[��㉄�w�⍳ߦ�
'�?Ƌw
��]��@����_�!ÁHC3[gq�H�C���.�ۯ�X(E(/Sl¯(:d�B�z!��V���r�qtZ��
\Kc�$�f� ��t�~ݟ�t�Z�{��*�L�����o��pജ�x� ������	|$��T�V<���bu���Z#zA4�!L���իQ݀�{�@k?D�]+��s��PO�+� =��Ἑ��/~v��<��t�4��$��E�d�].�\j�Ss�&��Q,X���`�H�?��7��Z��Z���SZl�l
�-8�©�dne��g�B���q��>O�R��D�l�pN�d�ZzEs!�W�#Vc���[^��q]��r�4S)����Ű(��K��SG�������|1&��
�CJ�M�^eD8zO���7�I�ݴhES�3���iր�l��9�����*��ab �L�_��	�@Q/U^sd#�p��-��֜S?�՜�Ĉ�T�&(��ټP�f۳ P�7ٛ��vPWQ&�ϕ�dʤ.-��1t�H�!(Ѷ�bs���w7���\����PI]�-�T`*K
�@G[�A`Qwg̈^���H�X� #��H��֐���� '��x�X��r7`p��t1�tB���8��5��#�kM,>��S��Ry�DNo�(�-f:wÄ�?Cf�v�grΖ�[�a�1d�����a�/� ��6["!�����K��uz	0�w҄�gҤ*�y���n6�(��6�N��3��h4��&-���0������$��z���<��ӭ�=E���23���A��96��ݼ�#�����߀t�R]s�^�Z*CF�,��P���RI����& �$�yy�ǿ�7Z��j!b:L˔��F�����%b$_h�����E�BTٺ�s�mU/í�lXbJ��y�e��ӈH1&'fK�Nes�������������f�h�-�C�L������������=��%��ܳ=�G�i{6�j�E���e^�g^.����cB:��M�ܠ�h���hϮ�?����H����8���H%��B��������wo�G�x��$6��<uңE���O������呪��p\�_�^������"�D"ݴ7�Eo���F��UԱ}�Q�x����]�QK���ㄿ�y�̌1u_�IjZ#뮡Ҁ�W� ���sV6�Y�\�]߮�>A=����u�59��q���Z�0WK�Y���O����}:*��h&����u���؜�e����]���vV��@�[ef�/Z,�G�~��.݁�y��T@`�j�"v�S?쉲ѝ�#� �3�h�X�[t�ټ�g��ȭ��m��{W��w�8��e���]K���)�\�e�z53��J�΁�-���G���x�rB���J�E���h�����<*��2�>���>J�5-U�xD�K@G�7�@�T�^֡fA
���wĝ~+"��O��\�@Q���՛�t��iLHm���j��x���e-��Z�@wK��\0U���;����~��i�]��-.��3��^?����0��#����/C#E�(���Qa0�A#�eɆ���Z�Y�\n�F��i��E��~�#�e�.��W�ܼ��Й��U���V���A�1U��W䖏}�*���xh��d;�3�4nfud 2�-�D������|�}������[N���>�ע��+U�������m�x�@I��\��p#i�NVC��0p$]28�Df� *  ^ ���_��Fzo��c=,'BM�4y�2ݝJT�#1�G<���6.��!N+�0y�{=�p�B
?Х,f�i�?������G�W�C�~_�d��s�ü/oKŜ2X�b��Oc���wr���Ç%�,�8�h1�z�RD�p9���d�^���3z!8�C�����9�}�v{sXL�_B�۶\E�sT�������9����*�����h�s<�v�k�t������"��
{���!��w��������3#�i�4�8�Y�2.�G�$\4��4�2����㚩iѢ��Zb:�W"D�ؘd��O�ߡ�O҂���v���IظY�%���z� ��]N�~9[�����1����4	7���]Q�`��H�r&���鵴�V�e�B�x�J��
�ۃ(����<����ZP�0��q�y�ۧ��.}0@ܧZpa{^�+�A��l,uR���EJ�iG�Gs�V�X��]�9$���hl_<�9l����hTU�*B��'�s��{�*ڦW#����آ�71�ͬ6(�+�'���n_A�A6� �W�!�����>2L�[�jo�7��zZ�R:{-A%=Y3�N�F_��*�-��0�׬K��=���pڡ���8kެ\I�?�*u��ռDg��˥��GP�h��4
2�\�fD��s�iv�ۆy��Dr��+V)��mK]��&�e���LT����XV}� ��Mrѯr]��D�q&�+_i$n���2	(����ę@�2k��O�JR]�� �D�����[H��8�0!�H�a�Ώ�ˑ�x�����*�;�u^K$�t| �AT�r�$(�*R�h���s�������M�O0��Z��bz������'R{�b�+f�{������ �ˋ�����ls���"��րxW���D�<.|g�O���|�T�H/�Y��6`|8=b}.?� 9��������U��|��"�j9E�j�I���ۡL.2.��K�']wV��|mNA��
�Вhw���C� ����տ�4�l�IuK�Ǚ7#^�ȍ\�MP��%���y���Z��̓� �n$��jD���s1�+����h��"���[��D�Z�Hz�Q��ـ�En� T   f ���_��F�����nY5*GF�3y�z
0xD�<�8�0�5HF�i~�$)ە��-���u�2wD��R"�Y��_%��H�o�oZ _v��~s״I�H�e�NM促�*O6}�>�� k=�y�3�2�=8A!Θš9��h9��קM��VЬF�a$��dt�(���d:2��He��9��K�/�eJ`���5�/�r���Ҋ���9��{��>��\M�:�2����}p��/r�M�ږ?���`���)RT��jsU��!\4�.��_}���w�~U�jУ̂|��<hZB�H���+��`#v��]��΀} �����=�hƁ�H�E#�h(��żO��zP�_}��w���+O������Zg�D�Zͭ�|W�ag��2Gü�o��b=#�����L�����$6H;e���0�1\�����G/�X����rC��©�������l���/�k��Vڧ݄�Х�b�)��Ͷ�$�Abf�0�������1�.�ԇRO���BLga`���[��I�-�bW�s�E�MGp\3��f�~e3�-�1
�\�}����w�,�7�^�آ��`�X� ��q
�:�����!�N�yC�Ly���.j+���P�O&v~��V/�1��
��ᕨ(lۉ@�DQ"`�����$q�,�5?�1��,�� ��/��{���\�����N����و�j"�6�<�3S=����Z�u��9R�|��1݀�����AF��a���\=z�HD9ja���Z�*@�Nt�-s�Mz[�r��,����O��,��&�K��9)�YN�=?L���k�kD<�_�GՖ8���Z^���Y������ gDpyk�a׫�5q�Ə�T�f�n�3���/���(�e2���e��8�M�c�h�#�jt��_���v���x��&�k��}t�<�[�i���P����_#� ��#y~����b�ӈ��qn:���iIf!�A�ͨ6�:�q��5K󩽢
��������٨�v^~�����4ȇ�I���0�A�[�ٛ�����㨕ω�6�홎����6�P|��b�UO��n-���K^Gy����?^*2�r����� nA��xp�����.�E��V�#_���q�G�f��L�����!Ba�Xf��:��	�＝�@�������I1;��cr���"�ؘ��"�[� 8�=j�5�SO��1�����5��?�@�IV]6��PkS�P��J�t���	Q���R���+Q5��M�'u츢@�G}u-1�>��\pj�-io"�A� ֛	��$P�X@���ظ�#�<���.�2T6��Dk"}��[i%+j��3v1� ��pt�Q}֑�x�Cρ �   � �&��F:0I�|I@Ȃ@�hH�/+tc�쿨|�$�|�;_�j;t���s:��ߊL�y'?;�b�r����/'>��3�t�
��Mj+,��A��@Lޝ#;ekQG�j�����H�uN#}B���ǥ`��^�Xǁ��[r��kũ��vZhDM�zV��N������f
 mA���8d�E�+m�ܺ+2��>8 ��K��
ɱ]����J�`���gz�c�|�ȄP�� A��ҩ��4,47�B5^�Y��Hл��'��:M�����ĥ;EX����� 1C��h���s��U�����V��i���#�%̸�ks�ti����I�N��^b�H��5��8x�f@8��!���_JIS ����q�*G?���ms�D)UyvI����<@�w��Z?�+A|��k�v� �6s��W |t;�۠��o����[-���L��.ٮ�rC��� ���`�4�vH.�r����vp2�Z�G����~3ͅ	�cp`�$~W��Wd_9"��4r�����(1��3#ˑ^2��C��_�mt�=`�#�tp��d��IQ(r��l<������l>DR'�;*�V��a:Hߣ��n��3��C��!ز�~�ġ�H>�vh%D�o�Ba�	)	�qL��.T����NB�n.T>���m��4{�ٚ��RJ�*
�JKB�'c�J[q�� �)�a�iv��#�	�����%�Ҭ�䈖:V�b�S �k�
�i�.�MMt�rTC��1�Ϯq��V���-��4+J�q�vzZ[�N���j&:�8�=���U�+�F��+\�:��e����&���t2}�y�+��9K{(�k���eKM��TG<���Ѷ��7%��3'�f�:I�g�&E��|]�
؊j�؛�v��n�!bz�r��W���U�$ӎTK\�E��ެ�V���[{��c��DˁУEQ�_����ǩ��!����&�n�[P� �CO �=�f�B�Wwhe1�Ks�/n��^i)RDBJ���/7�K�{�P���B����g+�
�4?���	��`�gu���Jk������B  %ġ�-�4�.�Ͼ�!	Lߡ�dP� `!��,��0��5 -� 
�h�"R��82�[(�|�9R� �� ����7C
�.y/uװ�*��:�kZ������#Qs�����ոW��|��
>΍���0�c�VO�p��	F0�2 
��y�� x%��'J���~��:��g�_r `   `!)��8��aS V 
 9���T�
�X���F�Ng�$|�	jan)}��=ן�G���q���&��C�[	⬺��L��D��]��Li!җ�X�ǒ\q|p���I-���n�ҀJ���a� �D�s~nx՘c�Z��)f�V�]3
�w�2Z�1ac�     !K�HAZ5(���pD�+ecF���S��MP��7����a�K9p��.$�R�%b�_�_���G5�W�[�����EJ����Sm1������&�o{{�7]�ٻ�Y��B\��T��y�a]�Ih��ƘJ�N}��$wG"(��g���Y���l��y���.���Wڇ�)�)�|�jV}������X$��}�S��    8!y�ҸfEQ�ˠ�ݴ�a��9���;�;�t:����r��tZZ��L��WfG�Bp��Oo:�[��mm�_�KF�D+
S�'8Z��d�,5ay�P��#�}��?���Ϝ���� .� @��Ś�9���E@�~U4˼;K�I-�Rl�Ӿ���~���GU} `     !���D��!X�h 5�L��BQ$�������m��J7�a��F�}��Tnnad��̭�v�����oC�"��~:r�,ө����{����`��;�X7|��m�.���,�Yw6$���$���6�n�����G�����|�    !����F
� �`E-�[aG�9�&30�6Ӟ�����6�snj���D���8� ؾ!����g�V�9�>��]�B����}i���^�Ki@R� ��������6�։�?0'a��f��v�ԩ+�m+.� �   �!�!�#�0�"(
��1�Ln
��*�`�@�&��R=-�^�ube���}C�&h����VAM�V�3�]��?`���;~������?o���D ��TDq YkI<!͍�@����ȇ���WFT"i�(���i%�qW_�wc�@f�(����M`�@�&���H��6�R�_gC��    �X��   �x����@c�32�c哴���.��W�^K��r�1I:_�G�椝�zC����=�ѽX���o=�8G����\����������a��䒼�]���޸�����>�o[\����\ȝ�[����Qb��n�k�Ō������?)��݊�%vl�U��X�{���g��^lgT�'s��N1��AS����c�HY�t��d3�[t(	�xֳ�ġ�9te�0L:=�/z>�LN"ܯ�A���rM����b�h�9�&��tW�M;����2g9�0���I.1�-� �Y�%�vQ�����QJ�+�<�.�[��O�W����R�@�z[��⫨�k� PO��R�u��v�b��o�o��4��yL��&�÷fg%*�"�W�?�h�!�s�����ls+��	(�턷���B6M�G�m��7j�R04ɲ��p�V�U�!��!7�N��-�	̥a[a��B��l��7�3��3<�6� ��Ͼ\�A������0�hm��C�eV��𷠗=ҥ�Uz=
G�b[�"8�"ƜI����tN���[!� g��3�Z����C����K�;�4︎q�{ld����� ╦ #ֿ�m��ͻZ�G��Ȓq+,`
X�ԓГ���t�iS,�ѥsb;�;�nDA�\�"�P��`ռp�,�jq����Z���(]�����X��@չΕզ��u�s
n�q����7m���e.ڮ���8�t��)��;0���p8��04$N*��6�B4�ww|�wQ"!,ov{��c�RI�����]�d|���V�e&p�z���h8/	�z�nD����uʋ��Z���^�:���pv:<+0c���-��z�\z��`�`�ђ��T��ODh+b��)׌�����U��m�C�\��b]�#�����a��v�OI�9��n8�1�X_V��
F+�]�9듐���4lL���gc�\w)���=�?XQo!���Zd<Y��Wji�Z��g؀�Uz�x�x��g�s���Z���?��	�YSpT�iI�6��gpw�૷4NC�#�g�c�aU���@'�?�e�k4x�����	�t��<�o���ʽ�O?��"�i�/^�ǘԠ:J�g�]�&�xW���E�0��X�5t:�5r]�ʜBR��H�����M2��Q*ė����y ��z-<N�q�Ap$	����ҥ 2Lk��sifこ* ;�2��#c,��]�p�VI��S7�B ����W˔��R[��	X��aU!B09���9�O�B�/�Z~��
��w��z���dw1��Q�Ɛ��z:������H���ij��C}�-J�$���u�33�0+��{��ⵎ���z�]J��秦þ�3	����=�q��6�*�^aV�>_��d`��Y��O-&�Q����^���n 9D"���I��e�0 }0�{�jASN�"�o��"*�
SE��tR�	��� F�\ָ��1�C�h*Q�{=����Ңd�2�ň*�8w����PWV\ߕz,��|%����g�������&���E���J�M�{��/���M��Y��Ý�q��!� ��u��1Qp�x-��N�����`���w��K�&?]|��<wu|��	�o�m:ˣ��nj-ҁ}��9ݖ�kw�o}\e���
�YW���x1���B�������yc����W���4����Ue��$o��5֟���0��f���S=�(ߊ�:rh��E�>,Mޯ��|���L�ĨX��cRE���7MA��/G�|�a���>� >��!��tܥ�[�>i"*&T*�O���Ə�gۚM?	����u�q���Ȝ��i�f���,�o4k3V9ъ��br@B<��d�LF�L�@FS��0����^�q$ %:z�GPюX���5[t�d�|b���x!�r����Rƛ�*0��
����y`�d�tZ_4�,.3��,��*f�i?:H	d�Ɋ�~6���N��5�~F���}B����g,�J����;pZ7�H�2��\A���R���@ �i%1��1RDB�R=4��ҕ!�d�oj~_l�t�YX=���)Qb��� >�觜j{���EO��s7�.c+�4Wă�f��"*�w�G�s�Ʊ��|�y8��J�-�3Q]��7hP�;�E�ul��0o���K�w}��4�N ��;������W�q��0aP�&�A�(=rE�~]N��n���8�ca0����4�Q4ZZ2� yvu�����,o�BPd�ԴO�I?���e �s����o^�C-ڝ� P�Ȋ�18�JEI:��6���Y/�<S�]4��ҫ`�+�� ��J��a](wA���B�j���L8TE���.;��y�x���<��'b������8!�p\a@Z\�dQ�hT~�۾]��$|�[54�54{�3BB���T�:ѥ��a�H.�G'q*.ID@��>�Uk
�i����8�W��JFĄ��S�pv(�G�?@��9��ː�96��iYl���^�>��I�@q�>����Vތ���~ɨh�u�AQ���9�ᾈ�T�2�d���ԭ����\78j�}s����m���I��&�֠�Na���"=����2�Տ��ݖz�6k{���˵�Ց���M]M� 6�"Z ����b�F>Ŵߘ>E���%w2Sp�@�wIg���a��mi#�_T��e�=	7o�~�}��9;n]���HZV�Z~_�3!�ܲ��,\Љ�:����ʕ�M>O^��麹�&�z<�����(|����-9�ܛ뻏1<�ފ�u��j��v��n��q?s��qᎉjNs��L�������0�16,9���)v��7���i0�W���+�|�>�&1��`@�g}5F���:�e�!�QsFx�a��8����\��C-E��Eh���2���\���汌5��#]���&����
F�2{E�d�S�I���������.ChO��;�9�:6�ͩ��@�U�]�Cx_�gI[a�]�t|���n&y�8zn��d鹨�z~5}�� �Mǡ*�P��������#�܇$)�����Tjߕ��L����vO}Q��Pz!@��D�	�T ��%��J�U���K�rD9�?.�n��_UBȫ&Ɍ�$�8�e� �� �~�m.����%U�^�$"�!�@Lbt&��9M|����q�^G��,�Fy�^\�n�w����kWx�:���oCVOTs��&7\��?U����	轖�i�M��U��\"%cG;�b{0��!�z��٤��d���L5�QG.PPC����i7{u7���P��T�2��+O
��n������FJ xv��9�%�n} ���}���#��t[��ۇ����v0;M٘ҭ�Et���C��F�#�i�?_�f4���?�x��������Ғ�x&i�h81����|r�a�6��T�-��c�o�����:4��R�EYR�7�z��k�j�B��&�f��B�3?��qX+B�y��X�AfJ�4DI���Cܒ�\�}�+�ؤ3s}<�|��^AJ3�Ԛ�-�����g� �)�z�n����2j[�4�.cqD�Т�L2R -��
6���v�t�ܿ�0P������W|ñ�����e�[�rbq2����>��Du��b����1I�ޭ�Z�S�y
�H ?�����ԞUޝ$�=W��N?��z�>iM���sv�>1dC����n�t-������:6{D�+e Q5l�=���nWP��y(�%Ƞ�G�?%I�`53Ux�Ǖ4�Ys�J_���*���&Q�~�àw'�YV���Y/����ћ����9�}R���7�n��i��R)5 ���Jd���W���kـC�~ԃmڐ�U���4�K��Yuʔi�TT,;���;�[G����!h���dJp{�H{��O��&g�|RS�4�O��@�vr./zx��X�>Y�a�Emq� 
�P��D�.|�Hax�,��K�o��#�����>���z����3K�p�*�hF���1_R軨ǻ3�KL7�ل�p�*���8��� ����n��FF����)"o��.�` U$p���X�ҍ:��W�%�P�Lq��Ui~<D�aqF��B�8s����<#��LH�� �w�A|P�������s䃟��7�24��~�G)FrL��!�|P�@�������h�i3�����[Q N���]$���ad�Qu�$��EX�O�,�x4�����������&ŀ���HP���>&@1`� E`S�M��H'���yO):���-񗲵~��k��&�.��&)iU�U���Bny�@�B]]pE�@�wM6���/6��5.�7{�,b�(�����G��68�F-zib[�n���!>�_ Ǒ��".R���Q,,��o������{�ހF�]�&�01��^_����ػ`������tM�$>9�u^��j~�����/�N�#�E�즄_�t��p�H�T�Tޓuξ7�/�vp��O>u�x��'�8cC��ZңM53���E����p�봕s�OQ��eR骈���Y^=y\]��	fY1jM6���Q`HD"��/�(���<}K-݋�Ȥ�e/�Q�S�}~�-��Rj̀b�����i�[Qt­-.��w�GވDv�hH��7�[� �uL�6]�LM�OEܵo�NM
Qf9^�(BM��uG�$]��)�M� p��];�ܔ��)Q_|0R�+�k$��;9�+!1��ꄅ\�0�m5QANU���w���@~���͟;E�[e��M�g�6���E�4�>�W_��u<���Q�6�#�ٟ�|�P��f�b*ڵ�!$�%�����d�3�*~�Wކ�d��A���+�AC��!I�us�Ox�"��9mm ��FT��]K�e���� ��ڝW �sU̕�Kc� �y����37�� ?�㖡p_�E@/�z��2�Nz0�-F*,$�_�K,96D/T���[te�vmnQ�d	��(A��2=D��}���,uRr�a�������������.����Sg�@�nRN?u<���W@���=c��v�y������{p�M�����2u��r?��>2 ��ٹ��3t���A��\~||�t��LC� �x�Ϣt$��Ŕ����O�ޱ�E��$���"�A\����_:�5��ץRo��̲��胆���c�J��O(;�	�G�����Nb�'�_7�fM������8w}̙*A�(:T6�W�'��)ac2�繡�^���Ϛ�W��_��ۥHRO�5���iX��%Z�8�#{�۟�w�*kcr�U!~> a>mRjL[U�|@XU�y��FO���M�[�nK����D\P����A��l�:K,DCo�
:C��3,�!r׈@}FU��[�������9&���5���N���ix��E�[�/X�g��U�����#���Y36�0e�&��Q������[����]<��S�K�d�7�}�����О;n������i������v��ণ*^c 2d�"֦u�K�&42���p��[\�3d�E�����6Ý`t���%���]����R?���j��U^�e��߫������Q�h,�:ųR�ͩ\Y&Ȑa���X�::�#���� ��7/*��
y'o�=�n��1���7�!7�@W�D8AT����mF�G�VP��������&3P�+TS]�o�Ͼr��������m�qO��֘|b,��!\x�lw]�/��9��aߎ/4�Ԭod��M���.M�,h��0�\��u����;�a�1�5cp��)gv�<���d*��m�p$�$#K";mfǘT�к�b\99��^A'༈��ߠO"��Z�����{�sπ�"A~�|���y����3�d�Z�T��3��{y<�צ�$�\���6��w�+DL�Ft���z��0��7�[B�=�o�^/֒�����!Y�e��ϫ���} K�J#@�%�Jt�����l!Ȗ|
�v��JK�HJ���*�	�P��zY8�����������ͯ/�̇(��t -p��\p�F�N  ���'W_q��~g��%�DR1��:A�v�(��$��m\���_� Gz:��
��|�Een�1K�U�<�N����NB"�z�������I��n��mO�G�f���B����1=24��
��/�5QH�S:n�̂��F��<����s2���/ �{�^1wOz2��z���&9�<������jƔ�ܻI8��j���h�t�V��9��_Y�c�����
����B�ڽ�NjS�~���m��0��O�ǜ�Jv1`D�q�koJa�it��%_Aq/xUZd��*�8p5c�K܏�_�א�y����P�|�t�d69���%�NL���p���\�5h