�����Jx�k�u�Yi�Y��(���̯���޾>�
4��T~&NnP�Ȭbv��z�#r��?��ZΜ^l�n'��Aa{_/� �yOP�xC:RgG��JĶ�z5�6��Qj�U晻��
E�O;W��ɵ����I��cv�%�
�^��o��d>�bJ���n=��3A�o�/'�uy?��F��h_�c��>�ձ&
1n,ϟB4)WL�����u\H�S��"���T�-6j?X��ΐ�%�5���`�/�]���V(�*���	!6͹���a��9!<��qc�Aʒ�ܧ-�G����������c/�}���軘+�P���������}5y)�ڟmd��3�f^��E�r_�	��|�K���>K�{)ᢤ��VZ	G˲�\s��8Yq,®,�~� j��D��h�}�pQ�]�pG�a,��|�3��N������˂��Ce�Uy��2�_��c�!��q#�}�l�f)�т5<��9�$��l��y�(`@I�1l�Y����6�S(�"<�A�oq��e���}l�mt���m�V4�?dԭ�d�ӝ<�*5LI��}J�e�)E+���V�![�����Za~�WNȺ��i�oO���lY9��T��o��i
��#W�g��M`�հ@
AQ���$߹�  �D�y   � �-W������"cƉ��A>�4�ݽo�Yl�'�q���7���j��1��pQ�b)S�� 3�|���+�k��i�<,�X|���@�٢N�^l�����t����ŉ���ѡ�'6~Mڳ`ܞ31�Z3����ܛBd�Yy��0�gX)���b���̓!e=�����@F,� ���Ց✟��2�\3��:+��1�M�q|Kvi�� �����N#wig/yP�L#n��|���g#0����eQ�������_X���XRk������>�1��!࿄���7F�=&T�M2�i�P� Q���O�t���� .� [�/�)�m$��q�{��^r/fXi�Z�h-����TCw9��ӎ�"p��'C�G�P�Ɖ�����kGLd�� �g碌�Z6�m�S^i^�	u���%���ί�s����G�#�\&������DK�O����}��R�Ğ޶���ϲ± 8MP�	�i%I�n-u ٫?G��� d��
��\FQ�2L%_�F��r���#H���.X�k�$áh�Iv
�����Y�	;Lu1%
i��QV$����og���p`"���b�3����`���N0�ލ{��.�V�I��}�݆o��X������bP�'-2�Z�c��W��L�TX0.$-V����6��J���HLos��iB]��Dy�����W
�@.	�{������z���U��:�ޤq�qSn�P���g������.s�R��� ���4����"����F:�h\���+3�3mB�$�����#�v3+o륕
h�t�m������M ��^�ւ*!�n]ױث�pq�J����X�u�wo� .�o��.���?��_v�;��Żb�)y�@EJmH�u�w�v��++����D��/�!��S�Wm��-�Oc�%