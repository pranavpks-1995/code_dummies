�bV
�hoh
/�@S��hY���T�Q��'�š���_X�q��~h�¹ x����M��� �R���$��kg Uf������x��{���`8F<��Ϛq�1!w�h�B����*нK$Z�!�R2�S�I
��f����c�Ȯ��Mv X������.6ç�iguz�0���j�ju={�B��r��:��H3��o)��o ��0`-��(�W [h�7KG^�#�Q�*��R��:�+�0IƧZ(��s[��R�*]�sr\钠�D?��vIbF6�KU�I��$��y��� vF��Ł��K�KݷwA�CjX�`�\^��T`�3��^C�e�H�oPp���%k-�As{�D���F��Y�E�ћ@�	ʱȱܜ�כ4���&�n��Q�g���b�z���y�n�T �����rT�$���|I��z �a��ǔ�xc.�6�դ����Q������-�v��i����fS�'��g�Ng�U^�V�k^'U��ղ4S7P�#��� ɗ�*C`�$���8F���U��(����B�ZoI��@�|L�����Z���,�묑
v�;����u�=��)֝q��M�l'������y��ЫB�H�&X���hy�I>�_c�	�����|��Z��JUZ�����(s��RrFS���<"s&xbX_�Jƻ
���c���[���a����RH�W�%%�~�}���c�F��"����3t��;+���ͧ]����T�