�ӹlV^���KcN�\���F��9!��L�q����@�ջ��ޥr��֭J���L�.A�y�T����6������5�q�e����n!y�.���8��K@[3ڛ���N���2�:*ҟgKJ��Z�z�k��;ncb�K���?�t��B��<�,�u>�R�eXϲʻ�J
��/�T���}�1b>�ټ�׿.��k@�Nox�j�9��-q9u6������ TL����ݓ*P���i���
R���.�]g�H��H2(����kΎ�ޫ�cy�����<�}W$gED��,�+�8{J`�3�(��qj���]M	�e/E���lقSC�ۭ����(@���E:�|Y�%Vx0yᷳ-� �f��J�����D���oDE8M4{6�y0*�b'M�Y��=Y��؍����@�J�ɂ�)�b�^WWh�m��H$�q�:�O2(�{Ԭn�s���kZ�H��G����ʞt|�ч�D��L0X�=������1c�Hg�ʁ3$j`�7�ј>t� �-n�[�:�;�b0_�?R�j�\P=�n� �IXb�N[��]����Z%�q�^�Ub��zM,ɗ/3E-[Y�c��9��,�#�����ભJ`�y��S���X�9��{����h��,�t�m�yWvH_X�@�L��m�{�niʠ�Hɧ�O���� �W��"q��m�EL���z����?qH��̯��z�}�q�Bh���k�p�]�&4e�~n���G1^Y��F���ѡ6b����6th�)^<12��~~3Ņ��ǽ�\U)G�.6ْ��}9��3\�~���F�2+��?>Q� c�P��d����{��tv����h?��k�Cr������ۙ+w/%���;=��DQ7�y�S��Hc�,�r�ze.�G��0��QD3��l��'�V��M�4��Twxy���;�>��P��A��Jf3k��ԝ"�j�4���aLTz��nFئ��s�c~8��D��x-h����4Е�{�����䒼r�g�[V1lD���َ�S����Jŀ���}V�<�`�_~�߱%r ��櫂5�X_~�H�l��B���
U;yו��A�6�*�`��u��O�+�(��Z�v�|a��̈́��!s� 0�]x�Hh�y{��Ե̣�X����{d�-�G�N��|�Y�D�[�a�N&#�t����j��*��x�=�s��%��*r���b�.�$��8�ݦ�SKz��[ަ��l7�>�g�*���hH��h�K��s����T�f�X�!��	Wd�So@^���B .��"���^�C/����a^��Tcv#Ӷ�>��P[��0q�F���!�� �HQ�Ng`��aa�� �ղ�4�v/�[&"X���Ba�׮|װ�L=t��;8��=�J8[QqE;XE)�
LZ��e"�&�`�?C_44!��k��ƚ��a���� R\��@��"Bnݺ޾	�S�:�[:��G&C�c����ʙ��H�z$;{z��P�Ӕ����� t3Fv�O"�ߧ��!Bgz�gAcX���Q���Ie3]��e;�U��F�v1sT��.K�"��g'�p��Om.�՜�RJ�6�g�V�����V�VcȺ�����S�lU�""��b����+��	�_zH�ޡ� ��H!|�� �=�k-�8 �{"����mf�1�ז_�rc=:��\X��C-qw����7����Հ��y�P��C��X+��bh��ȓL�={SW��u�a�;��k�\��:ڴO�P]5�
�N�O@Y�����"�~0!���+Z'OTm������Es�k{�0iR�yc�+���Č3I�������k�Uq)�x��b�Ť��C��  � �����,t`�y�ե���j~�Gkq:���`~�����2LI'�!F������������U��%����}��ZJ|�2HIv{��G�Du�Z#`�����gH���O��?� l����i,�����J����uE�.��VS��@���-��9���k[n�n��T�ٸ�vq��9᧐��khH�i��䞚fi�b�M�i��-c�H=�Q3+A�0���@���"<A��mxt\Kh<\+��N��qCW1;	1'��w�x��tP-_�g�w��6)�dў�����5D�BA��'��o#���V�B��37��U�"�$�l��h� _��=�Zu����F?�X��� ,6�,�N��ud�j�N~=E��qō%p��I�S{���Q
�4�$=*�?�08,b�ysIr��������Q�z��e� ��d���)�3�k�-���r}����#�<z��!`�:Q\ߛ�������,!���%�R��(�c�I+jĲ�.���\�&VM��r`�����B���� �;b��)���1&�׃��lC���yn$	�1���j�*m+����3���h@��&��htx�����xeNc�)���B�u(�<��4��*����Wc����P�v�o�`Z��h������+h\V���\�0��	zH��3!k�B*�*���}�z�(�)[)l��W��x�	zRf����³��X4"�9F:� 9W.6MW� �68^��e#����)�U&�T��Q	U����i䮷{�H2�Ke�؊����w8��S[�+#a�:���%��cʷ�ao�G����2�1�YM����(��s�d��?���_�T��������轄������j�����C�բ�l�&��`�����Vk������c�q�,�����0���>��kY��\kq�8���#ĝ;��I�B�r�S=[��pi?|�6M�'������#*k(�D�8   � ��-W���%�/����I���#x��j�Dk(	�4!�]�N��%�����r|,��T<�����$�I'��3b�:�ps-����ϞO˼��	vg�h2���Z�O���I���cT�) �'�@����c�xUp�(�柵���j���c�b�z���������Mk�I��p�^����>w\�:���f��*��^p�D/��ds�m*L���i]$	9�L���-DV4i��'����jL�(,{\0'��
l�(=�_4L�MJ�鰊�8Y��%0�w�r�΂vJ��Z�Z�?�*ǿ�ȥ����6k���#�,_�}T?��a��ϐ�2�1���g���E�̣���p�3�R5_n����|��q��|��Z�򀥳n�(i����9�����פ}酙b��q�<���g�r�Gɠ9x�[����v���k��+�.�#��t�h_K,�c����Hso`~>�:�.a�c��ה�w�N@f�+^�y�%�ylO�G�ԙ ^����ojSx
�Gm�#=��%�F��QQln$��?^���0)��ʩ�