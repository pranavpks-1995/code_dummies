M�<��j��3�g���okEb��������NpF-8*���~���'���
��U*�v�<nV� %Z�؆�r��f �g���$�Vּ�|�Bk2E^� $.\����K2rХ3����s�)~΢ѿ$z?�X�@zx�>K��?mtti�DM0'b?X@�Zch�n�w�>ƩL�AU{�=D�X�>'F������J�vy��t�_c�n�������|~\{q�S�ɂ?��n����g���G��p�q�	�����La���>�!�gQM�d�/�f�F��{A��¡o����3fcR�up��NQ�3�zU�*����r�d�<�tߔk����;~ *-�7K����S��������tM/�S[����B�P.�!L+��VRჾ����N3X�gj^�ljٝ~KڔcU�j��Z�>z73<�aI�D/|4���¥��g��(��r˱@|���ܬ��!��j��g��O�+Օ�i7J�-��X|�6ϖ�lh�XF���`�1�;�)��UL�v�o�'o �̿�v@�H�˩x��U�KOloW�O�oR��j�;N��?�V��![���OLk�M��� ���R\p�!�h�]�F�@�sH-܌J�H^tG�h�D�W*�ב,,M���U���Kn��b�S�ҏ#�=���	C� ���K���M�d�v��&�?F�~��Էr28���{�I�<C�x ��>5�,�ʻ����'��>���x�%��xq&`�
����W�.+�3d�4ۃ�K��[f<R复h��߬��C�m7�3*UH7(j��6���)\�咵�;֢L�y*�Z8�F��w  z �&�U� PM&�n�S����-	_?��u���a�1�	��Z.���{Zyr�J��H��(`8ߟ�	�4��Uտ�}�Z�
3����� ���w]���H��w�[���/�2�"p狿m��5�˖���&�^c1��H~;7��3`��pomf �A�|�Aȃ��z5�<�OVe$�����a�b1l��1��!j`��On 2g>:=�