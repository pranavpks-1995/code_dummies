���=�-�@�A���O�P�m<TPLS��7�)�a ��AnUqɄS������i�ͫثmY~ ؟�X�m�(qײ�2w���XH[\�]�2��Qԟ�_����:�?7~A����L�x��E!a�yb3!_���B�ap�?��n�߆Uj����ӽ@#�)�Q!P���'%.�B(o+K���Q�p	�'�@�~��,^#^�$F�/N�#��d���/{�����lp��s�i>\Bo��x�z�}ﷶ�{�S�jFf'�Yg3	F��@��#�~ҷ��l��쫓�]�x�V���&�?�1ԋ`T��s}:ᒬI$�q]h|yw��e�y��I,��K�ޒH;�2?�����%EQ ʭ�Y���cTxl򰹘�D�������T��){e�[hVo<^�!Y��
R�L�;�FV���h%|4�+l�@��F����S�툝��3��0ɼbT=�׊;�8	�LY'U֥��&�&I?ƺ�p|�Śnv�bF�XB�o�#W�%�E�rc��m�gH�wjlk2-9�  ;x����5G�EG����������!��`X0  1�]oo?�KE�˿6ZY"G�C�>q�:������_a�te�Mab�{/@��kVI�J��DpA�ؠ "�,�Ɓ���T�������tR�M�����-%�_��i�	�-�#���kɩD�:�9�"�����x&���U2�r�����2�� !��8�+�Pu�" �g�?\����u����HP���A5���ޔRaAz�؞��~��FksJ$��Pz�8�L�W�%HAPTrV� Am|K�6�ֈ,إ!�CT��%
���bj�9���	 �YݧΟ."��x�Y"��p�@F����.�J�`Q� !����x��4@%	]���w|��"EYeӜ�N�80���LՕ{��aV����qʒ��~Щ*�X*-8(�2G@�TX� Qf a�[.��p)���g��yH!���o(���V�[�2�H��K"�ibAE��
o�����6��h2�c��u�  �!�|��`&I��X���vD"C�{_��6��3��u��OR��k9�AII;�Άk�P��2��Т��ϑE�0��H�$ �# ��t�
發�r����Y��?��-G�q�X�j_)r����qrV	S
��s�Tߨ7�i��1T�h*��  0 p!��0n�Y�e%B�@  	�hjac4K,��O+�`��|�Zŷp����