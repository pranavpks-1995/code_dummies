 ��^y�w��D��vW47'4�k�<��Dz�Tǆ(�Jtv�"�����磥·�-,L��q�q��\zҲⅪm$zv�:�R�c���2P>�y7��Tp���(T����R��C�3c	�]�+f#x"��bA.�g�4�^ h���R����"��$-�Db +&7�\'lB��'���"�K��T�n_==���fך̾N��$F�<���Ř34NB�]? �����A�����-W37��<R��ޙo��
�_+����)���A�-���A�V2F�81�("��b\��H���>��Xu�E��[��)Ex��B���$~���!u��T�<���Q�  A�[�f����0����wP�e����3r	T��F��U�(����VL)F��{F��ۈqzߛ��P$8�ݤ]s��z+�2�>�â��L�n�Uco��s��I�IF�?iɺVg���Qu��^�)��*����|���#f�¦���<���v��^Idk���v���%��NB " �>zQ<�Y��oyy���>�uV_�fk��V�Sj��S�_έ���V"��j㧁�Z�oAB�I޼8��a����O�z�'�<�aZWj]�3BS�5 x����¦�#��U��S���Zr�QF�,�G���q�0|6c�=�C�����l ��E���&�'��Qٹ2U�D���� w\���,RK�sN���,�c>�A�\n�r���vK�Hә\{8@���m�����@`�K�J�]t]g�˶3k�P�Q#v��)����TKф�Է8İ!��rDC���l�&�=>��s�IL��z���Ё�$��B�MнrT���(��A+J�,ő�[@?-��B�Q��-���S�L�?w4�v3Jffe�J��v��ok����2X�º!���J��J������sz홃 bM���G�:����o��9Q+-�j
�tjʨ6�߿%P?Z�YH$��Ll�ר�r�]��V+{q��tss�pi�8
c�^T���a�3���*�T� �� � �z)�4{C#�4v">z�s�7[�l�,!�mpe�9�� .�j0ئE�+B��蹎T<K-r��l j�ܕ�}TazԠ;%��s���U���/�Z��𕽳1��|Z]O_`X�/W����^��KY��O� M`�&.'7�*�3�旳�����W�x6���B�ĔϢ�^Ubح�P��Z>��Յ@r[���h��d@�E�9�YsHPmԍF��U&�<p1� 7}OA�&�Pt!�Sf�'l�V1�@r��N/hh6���:m�7�y$��	�WU����7�����]�9]�>�J��+�aU�H:��bbG �r?1YG~���0�5��5���x:l	��k�7)���\n�,!)ٚh�\����ԁ�7�>�˧�:���ڽL��TI��3�x��:����\l�N���X���	�J"A��m��j궷K�=�;�wӕ���� �
X�I�Gi5��L�{W�r�3�u���P?�rw�'���?uI�F�3���8^6�2�=��Yzء�ƣ��uPQ�_:x(�jY�������?o�؉���Ӈ�����X�!<f��m)�%5�P�tK�8õ�v!f7t�2��
sLI�C �$�����j.���̃����.����;F���6�e��&lY�<wgTx�pB<|����iK	k\�)h��E����9�����D��54����ܬ,�zWB$���knG8�mpJ�i�.�ZOɩ��l���7��>�1��^��~ I{�N�k�l��Ӌʷξ�����7�&�4�J�R����&;~�ϧI��pm=�Hf8��J4��4SZ������kW�z�Prq�~SI:��/��-�4B��tf����I�>"@Sm�kc� #�* ��K�������/໯w��D�o�S�pQW�	>Up��N��R¼S�% �B�W����"��78��2qcN��n����rG67��:lJ?�؟��@�$���JF3�]���~����9r� 	A�i�����Ҙ1�P3��;esK��?��X�ѿ=j7۝�끂�s-�*��34����u����ڕ�f`ҙ-��.�'P�˰t�s�h���?����0J0z��obs���J�%�#�9��8��TC�-Y���k=0�<�'��9��p���ɩ�t�;F����T�kb�P��Ń;mӮ(	�?:r���=1���&��/��+aVĒy�2� �7N���G��[��5�6���h挸��p�Ąg��a8�����1x�1�1+M���,^����̘�5@[t4DS�
��N��Hއ����y�i$��<�7h�q?�ҿppH���3F��K'�>:e�C��zO����ȫxgH!�ucva��]�_-h���g�����y<��<�R�f���2��Х�k�C���U�qhf���_3���Ft�]���9G���r����V�*&o���٦�6�l\|N�W�c	���{̍�`�s�w��z@�-�3�3s�O'��?��F���#x=���2R=&�9l9�㫩���DO|V%��2ċ�U���x;Y?���ԙ�����A��L(:�l1�1j)I�!+�G���;R����@�bМ�\o!����K.k�И�Pi3�o�D4��x��nmi�f����o��bCk�6�n��,�,�>����.eݞ�'n&�xV"/�2!,z�2'�ȴ���R��f'p[ˡ����%�n�=t���>;���Rn5l�08�Z!z 3P�c'E��p�a~^QR�ko�a%�G��hq���ԙjL~��U�ݥ�|��q��N�e:w=�KК��Ʒ4k�Ca���Rvt�ֶ0A�ǿ3,4z��}x�u���J��C��)!Ҿ�%�ec�ɖ�����v(��)����s��V^�h_ ��A�����E�*v���]$�����I�^ঌ.����<ꌌ�A�{���W&P��Tq�lxM�?YY�2� 9ӏ��q74%x����#l=Mߥ�諢��(�=�+9����(��V��Ɏ��gLǃ� V�������t�촢��Z�z���2]��:4�d̂F���5�r��:~I�{z�D����	ß���B��M(g��v{e~G%��f����"��7����l�)=ֈ���10\��-|[�������(T�u1��>J+����Dv�H�W�Dfκ_�_���`���#�>J� �w��c�*�\ )��E��W�I�0�V��AaL��жa����	�6E�`e�&��"M�W��<,�@�_�@F)N@J#��4%@�vؼnD#C��L3���)� ����r21�M��!��9,�=���Cvq�k�qX�K:#��Q^ *�mYa4�ş�`��j0S�!���@��W��=�Ns98y�
?�*7��Θ�)�D��C�u�4["��z�nO�y�n�jS^Y��:y������`�
v��S�Aw֎�`
9�쟩�"\p��]`�"JT�ՕN�L����-Y�[������Q`[�Er�KK��C*>Kog��zތ�_� kT�c�0��:P1�
���Q��'PƐe�~�W$#�}�:��Z�N\o��o�c+���^ڿ�c�S2dÃki�]��x�,3_EJ3~G.�S�.�Y>��L9��  1�%RW�c�G�m�]��F��h�@�"�cئ3>�Hɲ+H�Nd�G��B
,�|��*[�'/��.�Xf�W��y0�
��MKhWa���>�&	Oq�8؍� �;#�l�!i�����eV���uf%ɂ��DL��k�~3�tU%���2�Eh��P8��Z.6�SK,5�eʮ��K��?��r;�K�z��B1��?�&=1V�#�~&�ݮ�7X��^V��ެ�ΙM�3 �ٖ�S�3GqX2˥�������҈ߵ�RK*�uD����`l�;n20���,7�����v7��y�E [o����6��	:ļ?ȩz�wpc��]Ȅ�ӧo���FHS!bp$R҇U��"��Br��)V�C��_���8W�b+(��}�H��U��1�P$L�P�8�u�l�p��KQ������g����rRyL�(��7�x7s�~��Zϔp<(�ѡ��[�8�t$���d��#jDxq� pk�4��}I(��"Di�.#��)�w[�,�Ev���f���#C��Z,���Ȩ�αf䱕Hr�Zj�s0��u'x\�����Q��V
��Ye|T�[��}��	�~f��[7_:MCHk�p��J,�r����_��bp�z�eϠ	���	{,�W���H��E�ȤV��:m�P��}���#��q��B�E���q���2s5���N��R�����i��ّ�Gd�&�N��}"�l��p��9��6i��=#3M˜�2\.�#�D%i�qu��(�xs^E{��|N1.P��Cr�iD��'G�Z�U�&�HH<뤫�_'�Aض��E��95a��X����ȟ�H�7�@��]e�mf�\f1���}�~�	�)�I���lz�s�ku-:;-!�d'Q�&+p���R���Uottz��׌��Y]�Fz������.y_ &�=�����V�_��`��ex4�ZE������ا�TS�Y�A)9�����ܶ��T�@�y�����(�J?�Qҩ��1��*/s����Xl�z�[��ڠ$q�-�Q�t�<��/(��سIM�is�+LZh��]O�n�����)�����l�K���Qs�+��G�9�]8d)���n������.nɟF�x��Rx{�A�V�P���G.�4��!HͶ�iw������A+�d�ؓ'��(}A�4}��Փ�֋q�׊!�`*��^)`҉%��ԇ刴�2�ಐ_A�@ļ
������w�a����kX����C?Hn��oV-�-
µ,^w?˧e���j�c�����ۣ~ӕ"<�&4s� �7ҽ;��{:��C&[%�saa�ؾJ&�����BƇ���;�	KNe�RvK�ɶT&���SՊ�cSO�f����t���=ե&pP��!m����yo���dx	\��u����SjNw�� :�V|N �>�C�򟫱��(��ٗ2!����<���]��y[sc����WLOorw�J
\�Ux=����g����m���㾐f�B� 6]�,zY@�r�\RZFq��5(���#ke�,�Yr�7��:�l 4D��������
���Bic�z_�����#O�{B�������z�D�� ���ߞ�l�#Ld���2H�����a�����a����ܡ��#_�)�s�H��+P*\h|�A�C�sKoD!b�=E���C1�r*���tr>k� �j��.�$��+d4�f�G�a���A��;�I�oc��.9�qU��X��,�����@߽�(~!�#�h	��H�U� ��p�v��<n����G]�!W�
��U�G��\T^�inQw��u�����#��-�!�F����:��?q܉D�t�B^)V�I 9#�u���m���DV;�, �n}�섰���2�C#_��O�@�,����/��u�24G��=����(�[�y��:B*�_>k]Ok	��Ӥ�9v�E�N��P����������%�{>>��h����Wot�����@��N�hMlё�4mޜ)���('|��Z(���#�	p�~���E&�00q����M�J�7 �ܕd�_��4�|8�(����i�9�>"FT��]��pE�p�2�YV"�q�\�%)�4�	�̑���L��Pz#��6<	f��<��@qVW�=���O5_�����qc�
��E9�����Wݵ�a��_�̽�Fn���('f��V>Om����nD��$�L"���Jp澌�cK��Rxu��gNw��@��4d�E�R<e�<v�����c���5CM�00j��Mc��A��n*�C���]Ťy�%���O��޾��*��~�y+�Z�ό�su@�ɧ �f��cS�&�3���Oɴ������`U�Qǲt�Ĺ��f�������B:SYTA4rx�M��+W� ���lpJ�`G�����x�m�@��	[�+"i���D�B*j�L�$'�F[V�=��
Yӡ@��#�8�|(�����w*��ϴ��T��;獳A�ҬH��i1�A���.^�:�3[0�[�Gvٖ_(v$�(UGo!�#(��I� v�
��3�$�����<g@�I����-,�+-њ��R&z��e����o��k����$.���c���/����&�Q�o��C������vu�x��� �����x&���"N[>|�6��ڛ�(-|\������IN����zw���_Ը�s�� 2]!�J���]@�/U%� ���e)s߸\ׁ�4M2\
�=��|͏�
����oNT��E�ց����,JƷ��`�/}���i�7V(k[& Nl�TҩY�{yiϺ���__���X$|�ej��mK\�DPt�� *I�@Y�M����v�=9Y���EQ�d=e)��4�$�_w�z8U�ݯ�e��\P&�����R�O)6��
� �n��������M��Dd�g�Hrf��Tc���]�� �u\�P8`!��+�t&����!%����ۙ��:��v�N�Η�O*���݃�G��nl��T����ri�MnC��%"q<V>Ny��(����@�`Ζ�C���,��.A��]<�Nv���&*��*�r{�s�Y��0��4L�ʽ�0,�\�Ea��  Y �f���,t`�#Z7,3
���� ����t}�"���7�Ks��٦�cH��=���輖u�ۇ��Uۂ7�8�)�CM�䧜Jm�G.�[@]�	�D�PH�fx�hb��6��^){�-�Sͼw��b��&��T�ݩ���?��41�h/�5�T�O�\��ST�k��vy�Ea�=;I�]��S�a�1(A�$vJP)+�1��<�W�n�{�F�Y���-�`X6�+��c�������I��阯#1��\s�2��1����v��;s�a���[?���d�]� ���?��․�$����r�<�|�52�s�I�����9���9�-�Mފ������m3����uo��1!W��
XO��\�<�(&g�ː� ��ޓ��#3����_�o�=M�r��"��>M	mV O��h�$�6�X|�e�&T�"���P=6�ڷ��I큮2��+Ċ��e�Xsb��D�Mj�K�1@��o�-��
�b"N��zaV��Zh�3�*=e��=F�1����?P*��*)��h#:ꡲ��4�����Xr�+e���B���"�8V)��%�ŏ���nˊ����"�*��N�W�c}<��K���<�a��&��Cd'^����g�}__��Ȍ���a��J�B��'w�d�1(�l��C�'#����K�pN�68h���Q;�}���Y�ᓌ
����%�n�)�e����MN�9���J�ˏ�y�o����C�`�7$�1\&�IP���Y�c�֤�'�PJ G��;ݳ��z�E���:f���Tʏ>�9:*5���L�6ڔ
¥3X��GX
�����4��ԟ��Ir���~#�K����������'�����y3:=*��Tdz-�@��`�O$Q4�K����F27d�����M�)y������ ���rkd��Z����w���Z��b�J��[1���i�|�4��![5��y�ʆj$��[�Cx��1Pkv�說mR2���G�?��g��|��������<�t��	�����Z�9|P� 9�q��حR�83̈́J|��$�Y�0�q ���E�Ǳ��H�8mH�̬R��u쓖��(���̯�'h�'3���
�$�#7�S@��^w%�^Qc�,�`=#����U��ޑ�����'r�� 1@y�IJ��!�]���Kj���<nH �h��D�C�'o
S��&q���~M��	m��^�n=�i��4���?C/U���������,;���pS/~���;HIh�Rf<+yuɾ���\ �K� h_��o#�뾊����G��Q7��o��	�
'ʠ.�v5��p �