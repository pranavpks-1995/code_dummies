ﹼ��Dz��]/���%�}xk����hek�g�������ǝ �H�]�]�\͈�O�i�>�B��ϩ�f�'������Z(�o`]�D`{�+ّ��y96!��e�M����o�� �&��*%�N�b��y�DƔ������}�\#�>��E�k����c���C����f6ʵ~��1]\RhW�c� 2�3�E-�޲oV�n��4�T��@�[��C=����9��	D��s\�𐧩���]��{xN^(����c�Dt�D¥�����c�	#Kq�[�u%_	�4S_#�{&�.�l�6U&y��%L��I4&�3�\�4�-Iu�$t��ǵ����D�T;#�`o��	����7ʜ�Cݔ44�L1����61(��o��ֺѤ�'UQ{�ɏ G�f�y6��9�	=��E��P�<҂���X�t�cE�m!S������(H����X�����JS:�'�O2(%z"��?&2wr�[���/y��/S��?�E���+Jn��G8*$�8Ա�x9$&-f���p�X(�K�E\��&$=K�c�Wb�Q-�}�qw��"�z���8p/�_cg;T�u��Q/w��Dd97=<���Z��G�3��0S�W�&�	�������,�%z:�|y΀#:m�[�¤��Mڧ2!�"�ٴ'GGˆ��3��-�p�t�|��%ˎX��[�)h����R�lO!��,&��O���(��߀L�Qܪ�q�| g��*7���(��I~z��e�^ȹ0�u�/�o.M�;ӳ-<W��	����Z���?�u ��_�P���q���~\dk�Ғb�ԤŹ�K��k�F�3Q)<5*(y���3�t9"�-� \�bO�dl��@EQ��9�Ю�y5x�M�C	���Y?��wZ�6��#j��s��� ��id0�}�����j�8��Ԭ Vj;���B+8y蚽-�%����5ߊ�V[`�$H���3�.4LQV�Y����Jyh���(��rg_����n�)�!�A���:�T�f3:����)VP��S�0��	ʢ�?7ۋ���xi��w8)#V��j�� Y�}��A�o3�HU�g�\n���o���>��}�IY��#
�o�|�-�w�a�S��&_H���8�k5	��ۀR��]�[u,��ް�Y�6��':s��3�+T�o�AyLі�BY
��U&����vW��*Oئ"P��"��J��=>Q�]Ǐ����-f��o����8h9Í<�0��T����2c����ń�2Tb����Z0�#@��U)��W��\����.d�R��k�����Ϻ~��`�Q��j���s�H#��~*}8p�{@���׷� Z ��9z�b���:j��ڒ�^�7w��L�\�܁ݸ�ӯ�Bv>ڽ�m�G!O�D���B�*�w����\DOM���5����2��iE�[ћ���$�-0���m�L͈�z���W�iY�8�&�#����7�g�5{���4�~��@��*E܃�Z9����j�	�iM��9􆔩WG��v���bѓ:�z8�u0��8F<�	�&X���r��[;�T`�oWv}�)u'
J`ۭ�v1D�D�]1,�*Cc���%������x�$�,%s"����L�����ȿ���F�Z`�o�9K<#S;�2j@��H,�M��^[�a�s�z ��	�1f���� �ب�x�Xb�-͔��Wk�*XNCo�Y3l��x'�7D�xoͲ�#�o�NKsCze�ǋ�2D�@�9EF�Z����# `9{��o���8:l)���]����igt]&�����6e��: ���%��o��`�7�|�c���ELH��VyUp��oVW,���j�70$&�5XL+�� #�����6NrU��c�K��ʂ_��P�,��sG������Ͻ4��u����Bj�y�
��W�8qlB�Rn�B��Dd�[�1��&,�Uf5���5�w�:���q+��s��+&��RG�]"���n%��ީܐ�ݏ��R��C`'�@�>�N{��_��󐄋#�l�;a�40۩�çR�H��Q&�h�֢[z	��%M�B�8~8G�B���Pʽ��>�\
J���DCת��^��HZ�~�:��&k�@MF�>�cք�u�/ZM��1-�E�u����+�&��ڦ"�* ]�h��2CDKR�Ap�S��QE��פ"��}(*/ې}�s������M�W��8�	� ���J���I�-�@��?���H�29�c�@>�!�K��ou]p@rܚ+�7E�=���/K�~w)�)F�lb�&����m���4��M�ɂ%8+ʇ�?�n�"�-�&�׈�
Chj�!��Lwo9&����dQW��E�y%kk�o��E�m��ˉ��E�
)�/`g��_v���