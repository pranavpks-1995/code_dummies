��.>V�l�B��VH��\&D���Jk��� �4 ��E�b�$-��}�OL�U ���[c}uj�1�L+.k�f����V��  !��!&HA@8���@ 	�?j�W�� �DW�u�^ �8.�Yh+�%��5I���z��Q�+�`4Ϣ���t�IH��ʓXM�d��1���)$��R�(j4�����Ձ���d�ۊ*$J�]� $��p1�
!� �c�e�HKQ�Q�?;U�Z�2cGi���ԆP�1�HURs5
�Pj���O��T   �Р�U��C��*]��B�p&��$�������XE�^/Uf*]gxx�	�r��:�yW3gJ�nuFlZ� �N��%l�#�`�s�kr�q��}��g���onh��긷/=
�sGQN����n��z�n�H�<I������Fti;(�t^.::�O�A�J����+�Y.���O�5S!w��ch[��X+�zU��������A�+�1�v����i&�:�YB�l�����g�L���3(=`�����������Ն���]�����[�}���G�3�&��"��3~�^����8Ӥ��b_.�V��)�Gfzis��o��B-ڋ���1�I�Ġq��C���Uz��'	��������`�[箉U`uh��/��rٚ����^��fhҤ�m|��dq��q���e�?��_��D�Ƕ2�r����݆��o~�9Y���v�r���||NT腤���$��6�x[���_>�L"� C��2ѷ	)��a�L����	z��aݗ	�S�G>k��<����p�j9���텶P(���R�^�I�(�+�����/k�R�8O�Gix��S?�ͫ�y����'d�<��H��]Q)��	z�nH#�6ǦaX�\��b5�@^�W��7>��qnƳ���V�"/Q;ܮ��C;gm�ѝ�|�`iٱŢ�-��@�ԏ&<|(S{����>��	�ID
�ea�L�CZ�>C�k��Y)[|J�����Eyi�2���	#�r߷[��!��N)
ڜy�p��p�;��g�X��浍aUU�_����^h39=��Ќ�|9��7/�����9�#�2J��4c�~-�q�P�z�MO�b��)�,�'��"�r�|�'^��9"�vD�I�|BUqaQ@�ܫ��'�9��+��}�0l�u�dժ�*+��bzb�}�E"��J)�XD��Z	�&\�����s��(��h�e�d�#Dꉁ�F���U�(z�_�qH���@ZkDX��7HF���qF)�����R��
���Mf`�^����2��U���td���^��}�����{��'�Iӊ�ڇYND��~�񵡝�18&�Z[�rg�\�[����d�-�I�:^�����Ǐt�.��s�4C�nӉB"_�C�mBO����U܎�r��m>��U� ;1h��oQn�I�R[M⟛���ѱ߽�y��ob�}�;OSf5ׁ5��+���EM���(�m䬯�~uӅ��Bd0�ߘe�k��*Ey)��Zvf�gX���w�5�C���?O�p೾�/H���BP�ӏ�a��|K���0�-�,:|)��;�K��KOT9�����W��[=CN/pK�Җ�)Q��8n	W�9���� NA��һ���vZ�ctP���0ו,Fn�����Ȩf���]	�CG뢂�dk�FCb���h�ayx����"�'7�Jh����Y�G�P�d7�da�'Y�j4HQBd���ɏ�\�'?uF
��g���2U�\%�H��?��Pzs�J]���yn�iGQ�n�r]���c6��=�3A��,1�:qۓ�X�4���Y Wo�qB*�Xȝ�Ήih���;[T��p�� =��)���Pu*���z �D5�u}���[df��\���nd�!��ZV��$�fG��w��`�e6�V��� �#��0�X@�Њ�osS$�?�xRqͶ߀n�"S�b�G�����JO)�doi+P�
Q;1�~9Ә�%���>p�r�ud�Hq�K# �"
ڌB�/�V\�2s|!����!=�t&ٲ��B�m���ʼn��$NE��:�C!�Չ=�tNǯ"�����:������~��eq�]�^�D�]a���z&��T&��"�;@��w��G`T��PJ��Ӈ�0��a�F�ݖ��[����|�v�