_Q0������6�j�\��O�ۣ5�ul�v�ѥ����O{)\�p�WHAq)ҧ��A(z��h���o�f�ʒ�տk�O�y�z'�k��;�.�q> �w���Je?�K�70��3�q�amϑ�J�PJ���a!�Xjck�
�c�fk"t�G`�4"@�SK)K8��t�Z/���v���z������w�W��
�k=��넯�o�#��CƎ��u[�O����pk�w��6۬�2��E�,�)!@��}W�\��m�7�+�?� +�0c[��`��S�
�=Q��\�B�3���,ѷ�k`0���e���a!v65U�@E]ͮ�5�N��[�p�J����Wr K����;��`E�Y2,U�δ;/}��f}���{*�F��'�r0_�!&fc�f|]v8���K�u¼�p	��gK��� pn/ 6?�7=΋���1Cӌ��[m��.n璬ߋt0�Y�F"��G?L	y���@Y(,�xX�T�E,�r뉬[��ܬ�0f��4�=f�;R뷺�X|�dɏ~GC�U�;�H� Rkݩ����K���k�79�A�K#�)٫��q]����̼^%f�����Kv��ӡL{��J|����Sa���Z/�s��*
'������%(���#^�Sȭ�).m�L��H�yѽk�`��yj���E�]5׉h-3n�Gk~���]6E��	�,Ke8V� X�h�s�� �* �!�]u3��|K��n����0.j�o�d@�����ޢ�D��b!�S���ӭ�_�=�
�s�H�v��Il�����G�P���� '1�IPd
|�#>��^�g[��{H�eNH�aA���]��~�YrYC���mN2G7�u	(o��xk�=9�������[�7�iY>3�G��KƋk��h���Z�Yy���H1�2�N�(��g,@ǒ/�	\����V8�e��M�