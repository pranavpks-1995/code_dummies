package INITIALIZING_THE_RECEIVER;
	module program (Empty);
	endmodule
endpackage