BBn�/S"!��j�5j��g�ef1�Yhhȵ��
�q���;�O���4��\�![�|�3��^g��C=�d�
3�`�b��ƌ �M�Y~����&����Dd�2�>�"<�T>�g�k�s%��h��~��zј��pM�������Ԑ�,>�V�t8��`�F&TTǸ�*������-��4@Q��'���������g#���L1�B :Kp����䦙��q�E�a�
~���_ӗ���?��4��r�d\�8��l�)�-+{��_�&R�o�f��E�9������-�ثf]%�j���߆��{��
'n�M���+�����[�<��G|س�J�w#ac�P_��"��c;3�qw�D�iGL%�%"������G9M0�(�?FF!���Ʈ��6�����w7�,+�u7�"����	Hȓ|��/E(4�2�ŏ>�1Ï�.M||쏵G���h��z�>	��h$��葑��"j ��w"$������DڗhE��9F[���Q<�����N¸�7�*Pm5m�&H>�(T��-C?�Q^�J���Y^���V��Th�^��=|I�����p��D����U#Q��~�i�II_�P����-m�m5S�ܴ�`����n������yq8��nV䛚��[�
>B���$�;�Ki���=xwfn� �U�};�U��bjR��+�e$@k���}&���)��,�ox�v��r���?8����-_p=��nc���87�vH�/��t�2�����6x��T��&6Q}uݪ@����zb3����#�0�
&��W�4{��V�vJꨗ���mvq0-���k�)�}
Ar�+ݬ'�s�z����=�(�ݏ�s�M��-~���\�+�	U�{�C�&�V�v�v�qoۣ�fHL譻�Dz��ݑ1�+��s4x��4x^n�����uk����� o׸�g���{慡/�cw��kG���a����V^!�G������__�"p�̴�|�O;��0^�(Rl9��nBAM�xW#wpvi�c�k�X�E�	@s/�x�͔�_�j!m�=�G-ҝM\3��~y��C��!N�Է^J�F'�ޱ����&���SPU���cV�'��9
�����z�o�hH��������\�+��D�#�y
L�3����X7.�O�*V|V#����W_ǅ¶��Ύ(�)���]�#FQ_��y��N%ʕB_p�<�`�,����l!
�A��rr��8�Bm�)�Z�՜L�z#�(�6��πD��#(��
6�!�U�E�Muʶ�Ƈf��'F>B����H���_E%D*Xi��'m�JK�)�7��S39{Qc�<�~(�?�C��XY [�km�	J����@�y���q�;v�����MS']�
�� ySi�H�;���G)?�D�F3��K|�+�ˢ�)C���ᖧϕ��L�=�WJ|T�ӃC�`s(�ʯq���L�0��漝(wY�6��"���0q��W�/�2��7(�h{�;��n��{�K��C��h�Sid�C��a�G"JZ����4!)��d�zf�f��weޣC|�A?���W>�ͪ���$�qѤQ���a`'��:�ϗ�A�v��"8�x��$I��)i��L%Nڑ���M�vR�K\�1"�"��gi2Յ�ݯ�� u>�y7�v�W��x>i*p��qg ǭ�>6���8�,J��h%�U��}3��f%�r�`i����Vt���)P�ה&0J�*��$g֘i��WE��҅��⨔ c�����.KR����ť��,m�{x65�j����b`p���)/!w��0x�����df}��降Ѿ�t-�Yh.�c��F>Co��ǰ���:*I