fP��8`� G�+��Y,C�Fx�k�d��������E�
I;B<F+��e�4s�� U�?�)��C�4� �̉U��A;г��^�P�gñ;\W���!'+
�I����Os��k@Q�5�/���#AΑ���o���Ѻ�-��PAF��s��H67��[R�%u�%�y>�Oأ#\_�5�⹕gW <�*&c,�j#o�]=�LJx��_T�]�@$���*;�s�r�e�A'�1�N:��~�ƙ8��[f&����8L��pMג�h������eI����I��� <�3�c,�w�س�70�15=��O��O�����`�,�|��a�ȕZ�_q�F���,9@5��K`���x��d��B=C�o#;�H�a����4i��F}-v]$W'i#�qq��2�򇻾'�?�ҫ��$01����o��	w"�����#T���ʪt��'r�����$MH���a�=V�����=]K��]Nѕ]!�rM�,�)RW
�!���{mB�(�H/U�D���[R����R' ���50��+�q�Do���w��az�J�d���:Br]#8�q�u:n���g��S��pT)��TRi�=̹Q�	N0 dE����[�-((�lz��u��c�+�ױf�x��[��
p�ل��׏7-�hV�]�9�49�%�q��9�m�$,�\9�j7.�@���)���up�'I;��a,�6n���7^ClOs11Ty���1�*�,]��֣��I�;�7�\�q(�7�,��07̃y��eJ�yy��ڙ �A(yQ	�m�g!�L�6kў���:�xEͱ�ӂפP�K_�3���+h�����.J�=�t� � �E�
�  � ���U�$
�d�ZV�<@��9Nlt���@c�B��ˤ���J�l��|d�e'�fz�i�&��k4�X�;���.�����HwZ�fO��V�`.e���qA�+]u�\6�jτ�s� ��psi��d�� n�]  �s�b�I
��U��'��̲YJp�'���Y.�]�T�������,dX�ܣB�0��@��QX~Ȱ�H<����(����O\ބ��(�,Xa�&w'����;�ҵn���4��{�rӥr{��~w�I��3��n��O<��r��c8�嬓��-���z��vm�ć����;�$Y��e%}S�N��칻����tV�L^Y_�h�	EH)v����k�(����mp��j0�Ƹ���O�ΡZ:�yXD �FV3��1-]3k��ki̲�� i���[����p,�s�(:�0��}���V`�����zF�cR�^w�B<X͸�/B�F�Tk�eS�S�2�atgi��CI�X�V;�e����MЗ#A���;��#<���ڵo&��vB��͉ ���Z�۳S��-����.DA����h�a��J2v3[��_JE�|�ߺ �Bݰ]��ׂ��;|�m�L��J��0o�n��L��"P�c�M��	η?���őn�P�
GYf���E�L	�oJ9����	-��=�F ;��?�|����9��&xm�"��׮�%ZI�)k|~k��S�g�&�=�{d���Z��>��;���8�+dl�[�mu�\�22m��H�����9�[)�W�5�Z� b��Ys��o��ŋ|/ޓQ"�=�g��UU���Z��������&�EcvEY/�3_䞤�W �i�h�<Bnx�L�(�.`�|"�s�����ρ;��u%0�4��e͏����w��&~�T�v��U�P��r�-�m��{�i�`�=���f���w�v���z\3��fX���g�V�@pYX�O��9��x�	�t9�M���n�.m��܏��'V:�-�Tf���z��R1�H����k�����o2-iC���D
x�A��6�!5�uHp��&��!c��&3`	).����)g%��E�~������:��!�$�y�G���|��O�������b��,��ºx�V��C�D�<{A�2��(R��V�$�p�~Y/�ۿ:���Т��m�jH&ga̲�غ��^����ǜ�Pc[����e�yl@��r��90ܘ���ǔu��R_V�9���{�j[���'�ci|��@;������7u6q�%�{.�jҬ�t��R ަ��Ta�ɥ�#�b\�%��(3�L.̄v+�o��|If~�i��hOk��+�ܬ�����,O��6��Ɍ�߉���Sa��>x;��;!�1�x���֔3C�=�͏e[hQ�g��9+��E��:꓈��T�-5��������_��UGx`k����k<�,��t">;�~��G6�PON�e�)0�쟘���WK��F��
�   y ���u�$ �Nkԝn؞+�6�ߠ�CD��PoC��#b�����'+<B�-��CX@ `y�td�OX��څ�.��q���&a��ˆ��S:����Y[lN78E�q5~�P�u5��;���d_�v��I�}Z��p�\�OKΫ\�rD	<I���.�v���t�#�Ğ|&��S��P���Gh̒�d��f�F�I�az�#ֻbNOd�@>�iɃ^�>p����kF9�(�:j"HX���'Vy��j��}�5��?���}9ܪ�K��O2=�R`m
@	ꐘ[˘^� n�_� ���a'����l[yE`z��T��`���l@̜��GO��CS��:3Mx��p7r�Ӡ��
:���ݔ,8��L�+����b�@?G�GF�1��n�����	0�8mf��'�N}p �UUF�����Ҁ�G�`�x���
�h���W����'�R��rxk	�
��d}pؼ���sT�q��
���d�W-�4�'��
�#����\/�k8S�<l��S��b;7S?Vv�]�-$��X�-/\2̸���sTp-��	� �'�ͭ�R�yXb�(A�Bf�wh����/v���.k`G�SP��Ӊ���-F^Ըǲ����'x���6�ܥ+�����K��Ҵˌ�F�p'V�ȁ8w�N�8�U��|�+P���=��Ltʐ�HO���۠kT�$3W�⽄���r��x���zt��1l�@3��_�����`�N�I�Jg\�T��^���<��+@ã�}��a[#H�$Y�N�[`��A��K�d�bp��İ���B���4�eի�0;.�����A\L���#W3G�K�5Ov�1��w�$�%R���N��G� �e|��
nn������3�Sѡ�%���K�"���u���.`*fV'V�<胠-��o:HO_��Ү�/xf�	��޿��8���.���۽��[z:&q�_�H�٫ ����G��X�7�沫��I�;���ܖ�}���m���p9��X2��Q걞+���WgR��4a��&Fu���K �&_&`���y~(�fÇ�͙G6D�LVݡ���D� �����!���9C7M��60��tA� �H��"ȱ\v/3)���#�9�M�	�1�x���A��ތ�Lf�Te����6 Od<k}v�M��p�P)y{�A;�T���ɥ3�N������G\sU���;� �[�he}�I�O���"�.xv ���\ |:�)�-��<�<7m_9�X�א���)�q���+˒�g�!GKP��)��ީ6��W�;��n����,}�3,�9�o>��l�z�����? �=�Z��sXn��R,��;-e����T�:<pza�=>9��hd�,3$�Lk���J��;Lމ�Q�d>�횖�3;Ð \�C�Q����	��~L����SrE�n?����]�9V�A�3z��kˆ�HO�ݔ�`�K"������fU���V#e�����EQ\���'d�:��XG�+^��3��%�h�z�k�k@�/�25j"��h1���ǉs��Ȇ栤�! �F����+���:B� lzh� �9v,}yu�f����������vNr�z��L�l	'1�T�E�    �"-���� �h��SJ��3��_5��3|K�yP}�:@�)@�&':@�����v�	���C�B �n8F\�&��Lk�;qĀ�G��{l��?�����<1y��t�r>������9���N4�`��*p�<B��Gv�����r��C����0�a�:��x@
��C��AK��:�� ޜ�%i�S� >�ü�� �c��U�ے��`I�.���Dh
���r��A��,1�>*�YO��I�`��l��h��X�i��M�ڭ�Z���%0����d.g�OaT�c���Ur-
��`B<}��Da������O-�C�{8Kn<��A�T���d3[�r����<�a"�[%�)�Gq^�iΡ/�4�x�w@i�Z5޾&��=��Fn��B�-��o���wP*�~�U!��MG/�,�Kw����#'���/���5<���[aF�V����qXا�2���{w�\	��L`/x���H�Y#�H�ҲӔ��L�K�6��,�Ff9�q1���/	�ɛ�Ia��F��,)��{����Q��sr�z���v<���HC#��A�����4�ht�[ڟ1�� �j-�G����v�@�o���9u�������S�ȵ�3�Gǿ��z&��v�~�S�����5YWz��f�̦F,P��H}���pFs�>��\r�{	��;��[�����x	�*0gI�u��%!b�J��aʳ�ލ���_ܟE�2OɐO�~!�??�?� �S��3�a@^���N=�g aJ���r��h����J�`���G'��h��{�%�:�{��W�{���j^%���9�B��t&��>�h]I�,���S����95��V[�}c~��ty�W�+�Q����XJ�)�?��q�bO��*$A�=�"�<j
�w����%K�D��EjJ%^~�˲��I�`��e��$�7�1��d��Q6'
����n�����]�)s�6��/(�����in�M95o�;�*V�ƹ��Z"v�0�o��>W��P�%�e��a-�����&�}G'M�
8KA��n�&νTs=0a�¦��7ϑF��:d�9j���m��\��Ä��a��k��,��#�P:[��k�9Un�eL�- �
~�,�-V��b��� `X�J5k��8�J`:3�a�3i�ۊ�8��^�V��9��T/��4�;y��؟��ԇ�Nj�H&f)e�!:J˄Ƅv���/8�w���PB���쀣N���   �Ѱ�U��C��.Y�1R\����@`������ ӫ��*ˢ��ћʑw�j	Q렅XK��=��h��,?i�~���m�iK��Pif�Վ�U���z���=P<�];<K����L�?����A��p	��{��R��n5��jP�w���FNR��tҾ��;��n�XU�j8��t[�Fݍz�c>_{��0@t��;�?~)B%�R�5\c��h
����������z�yfb���'�6=��'�'R*K�'�L Ч[��8~�?�|