�	�`�Y���������x�6�?���#�$Y3�P7q��0���r�rr�^(�%�.��ot�i�O�����jDcp8YVG��!�j��=S��F�I���4�3^��?bO�IE4��#Q��%������:�����m�D�A�2W��K'�H�!�c+$Lu��D��i�0�4�;;�� �G�8_ߘX�0Aõj�~Q�Ϭ8�;��HgټoX/C�$���x;��,����}��[�� {��t�}^|�}�Lo�G�!R�XM6G���X��ΞK��/*�R[�h5C���.���������K��&e��Dn�Vhog�GZ��DTt�����TueU�++��)�t�R3P�;�^e$���#9�J��z��潥a�#�/�G1��@�ã��(=�Mil�q� H�K������Z�	8�vn�1:��ʍPr0��9�:p��{[%��=l-Ox+q����#�t�kf�.���K1)K}3�JPٻTi	a��-�&�= >H$f]�1������6��p�)�#�^|kYo<�"�cKq�Xv�Իr0yr��TJ�J��zo.y ��� �;}�1x\�H��	U6�T�dC��5ur+��~Cl��q7�ZI��.RP��,�ԫ�~掲����^ܖ��"��_� �`���=��TCۈHb��>�>�U�i_W6�Aq6#��4�qas�E�g�\	�wV�#���Vnģ�H��^�H���b���O�Y���jA�](������M�Z%������wq��W>(S�ð��~��D��S]����:� ��.~���|M㲻w�jwc�.�e��3��>�DE;��ĉ��p��ﶕ	`j������uh���Z�z<&�7{���ԭ,������ee������*�@߲!JE�Me�s�h׬�S�pl��k���Xr�*��i��Uq��@?1���8]�쨖P�ui���)N8e�ЙV��B�Hg,���<����Q�N��^k�lZ���-�o��F�vտ�Q��=�y{���D�p�ݍC�O_�#��ɍ��i>w0fݧ"�}�|f�[[�ܝGлG���O�!Q�o���T���k�^Z���h�*�1<?�"5�X� �Չ���J�Ś��rN\�����6u�O�DՂ�L��՝r�u��D���s֨��������X�x�ɭ\�,�|�W��-�O��Ǚ�)2R�<Y���R��ڣ!)�j~����y��%gs��³�0�8�e��|4���@q
,ZfK�ˇ,R������q���A��,���O]����_�x,T�Y��P1�8�