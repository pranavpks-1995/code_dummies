>(����Q���iK�AJ�k�4Ӿ�P9��X�]�\p5��w���ڿ�*��#`���AF�Y�S�[Vߊo
m�q�-<ț](
ƙ]�9���E���;��o����w#��F�8��@��h7D�(��0��<�V�[D�ғ�g�{2�J,��3-�;{~�z6�My��Ļd�Ս�,Z@����=A8�(q�ƽ	gk���ZѠ�Ek2�ڸ6�6���y�� X+G����3����BU��   M �&�u�zO��B���ƌ��ÅF�j�o��*0/�7q��j��~.r]/.��hy�8��!tW��{{�\���}a�w �j�p����^a����Ch�D8e1�	`V���N8��Ï�3�8�=���Hx����.�8�fCW�n�NBAYM�d����m���"��NT7����@]5�=�
�b"�L����$��K�w�O��cx�f�P��FSd��*fԙ��Մ�K7����v��ۋ�X��a�C��2���P�����9���ho(�����GUW�ux`56!ڐ�R���:��l�{�{t"��t�5�l/�W�.I/�Ǹ����G�*:�����Wr��Js�П��e���
�	���9��@���m0��b 13��y���Sɨ������J�0����0~%V�u��pu�mi�JZ�J5[�U��;-f�Uĥ��k������,�
j�;�\&��@{��9��{�J'��?�+6���o���ı�!�5����������z�	�Z ��L�{Ӆ�}�\�y�J�Sa#���'o���Ϛˌ�+$&D��v����A�0(���*�+ �Aǁ   � �b-�����\�i��<J壉�:LV�k�[%��
jix=�o�3�0f�-87�!��� �^�X�5`!V"�x]�Ä�B������B%d�Ǳ���sqd��}��o�3I�������q���=z\nM�$Lo
���s�ơ]�(��ҮE%4H�y|���v��G^,~����t�}Lgv�3�܀x��TF{1���:?�00d=شvbgz�hc��a�dq��7�ZQB����W�;ts���gc0�-u�Gs؀�a��sCY)sʍk�h�6��������ԥ�ޔ������&�W���}$�{�c��(�Z��X�����ҾV$���W��IopA,h֪F�+@Y(�Xw)�z+wZ��O���W$��r9�Ҽ��Ac楹j��&[^YE����f<۞�kF%jo����\�~tCᒎ��d��~�2���(�k�4�Xw����#������ They thought Joey was a child?��~�E���������!�����el��
A�:�`��䚾BF5��>��Q�t�������~= wM{ȈO��ֺ��z�Β�;�4�7�R鋐�͜�-d�
*� �� ���o�(�u���d����|�;A�`ыlnp��J	 m�T���.^ �X �!�� ��D	d1"�<W"��R�4 �D��<�{��:�<*��"`��ٓT�P�������;�|s<!�����B��<.��O]8�s�������h=WN�ܐA��?�� �Z�� A)����q֣s>���Dn�1�Aϡ�5w�x^�rj� l�V+5"d  �!��`H�!�F�WdQW�� 0�Dƥ"�kH��	�4t��w�р^2�-�}0����{��%���w� �sB����IqMUE���gߺ���3K�-�S��J�2����Bxf:� �d@bh {� B�l��{�6��;���!�����!UN��kmA�  !��`\��s�@k`�u`3�>^��s47`B�����'��� ����z�$�%�Fn䄔-D��8���!-�X�rv��h+:x�Či��&@B ����%wt6�V���Ey05.�2���z$,  ��^���*�� !��1���Y�6; �WcKh�Y	ܛ�{�֕-U�ߓ�0����t�.%&�'��Mq�)�bXM�3ܪ���.��*�-��YG�n��1QQk�.@�u��� Q J��cK���p#��u�Cm9��!+��Ԗ��?�R�k����a)_�q�p� ۤ*���Z��� �!������۪�5�`:j��QA]���ʤ�"�:����T#�ix< ��P���������8��G� s���]�T/"|L�� �E�V,9c�AƁ�()E]A�����P3\��i2�UN
C9��V�(����o��  !��`ܵ�۹x��x�`-m *@�1�4�m�	��J�f8�f�XojBW�$DCS�����F�)�fH�TGGs�-�)�فmyp!%gʿg���j�hB)H�Ԙ	�H`��H�QV}�'��u0�m!7ZVf�}�5�U6Nr<�b�J�ɂ  !����p/��U�`*����&"�?��oi�E��Gul�Mu�F�*��B�O]+�bL��{��\� DR�s]>�i�}��Z���2�mg*����v��~��f/ &� �8B@#����w�М��+�o�ڒB(����TCߨN��6=�#��T �P�   ��H����C����|�1\G=\zE��BSe,n^�KG�0�xIoy�'��@�ȮIq���\�u�'x�n[*�Q���(�LV+�����4<�p̿�r3�^=�O7
�=�i"�����9|���&V���$-�Vq���W�KG&
Ϫ�:*rM�2l^���}RqOWYSp�;)~huEjڹ���"�i�	�4{��z��#V݃�+r�X)�	TP3��)>Z�e9P�$%���2Ys��Z����<��qV�Y��2(֟�r��z ��m���?�h�{+݃�N���_���1e���V����Ϗ��tg���	ۜ���~_�Q΅�~S����&R�lE�Ϩ��?ړ�t��(�2:W{<X�<��Ѯ�d�ܞVk�U�"��V3x�C;K��$��̘kS������k�n��D�m����__���;��a�6��;��1/G&8.yq�)�օ�����S�@z�y�L@orW�I�_�3߀Oj�v���dQ�
+g]y@�=��Z,~�>e����u����pmK�
�/8�g� XU�Pv�菹f�%���t�-/T�$v9���v�#[�}Š
��+��gQq�!�y5a;]��W2��ѥ]���ڜɶ�^���-�!7���}��]y���NtE�]�a�=9{~�i�:�{'1"���8��L��8P�!� �\�|˗\S�����U�=�v�gZT��wN�M���qā�~���3���s��i�R�a6�g�݅��g�����e/���1�45�47�J��V�H��џ���3]����oA=t��b`���p(�fE;�IL��Xepy�<|NU�X����AM���
'�m� |�P "u>26����!���Ұ�Ȥ�k{�/�4�r�2'�B>F/��ʻ���A-]a+J��PKO��YxI�(�U	�>#�D��Gp���:�\R�i,��g�2v��e�b�h�j���;c���B�.�D���`�WBw�F����KD��*��n�ZU��=f\2�̥uK�YSj�g������|d�F�A� !���^h1v
�yd��E��*�є��*�{�v��2�
`&2TaM{���dW̥yu��\L5��K�4<.ϹN��?�	����O>/p��-7��IE?[Օ�qt[��'E|�ܷ�i�̶q7M5h�U+��B���s��"J��o���"�"���+��蛀�VXM�Z�I�5�!u:���Tv���$�bП;\c�[��N��69�@�
�7RZ�AF4XO�b�Ŋ΂��_��h��Nf�q��KՐ�/	�{Wvk