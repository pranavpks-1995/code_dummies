9gV5SP����2PMڿ����?r�(��ͤ�G���k�zO��"D�3��gx�0g/o=��	�{�����&�ˍ��������>�J�t�Y� ��?��8�'��{c�8UlQE��矄G����y���F$��n��,�z$��"��~R��f�R�I�S��A����U�A�i@��r�,Ef�<L��3�:)|������;�\�wd*R<ќÙ����o9/S����e�E�h��Ɗ��� ;Gϲ��g�Q��x3�dc��aã:���"� �0G��O�/�7��V��+�7��W�`M�f�����d���<^�y#�'x������ō�%��hW�e^�e��n�+}���9Da��&��b@��C_�5��A�z�Y029�DR�y�*G���P	HRNHѳ|C�^�I�]��VJ�,,�\uJ\�sn�@p�$�6�R]oԔW�!3#9��~QY�E�7� �ץ�d5Cp��n�x�5�0H�!��V=�"�]z� ���	���R�۳NU�h!������<P/_�u	�J�ZP�z�̊�su��֏�.���}a9"����*I��x��A7t-����k���2b� ���wI��6�WM�H�w�9]V�%蠀�ů�r�RO%l��y����t�d�*�+�5V�*���0	U����@�*���\v��t�ӂ�5�/]��%-W�z��+�R�����^�������X2{6���~�X4��q���@�6�9A�/l[~