��Q����L��:�^��;���5r))�h�I�!t/�$�����kMD�J�v�n��v(����],-�1�_ǔ�O�<�A�UQ�	C9�{骩�)���&���r��&�� e�C[��Nu������fe�ɞE��j��DS����>�g�h+��9�xla՚�3��"ڽ�6H5��{*' �6K,�����aըY�Idy���؇.��P.`f3ߌ��a`[.)CW�v�~7�Ⱥ ����5�	kMтs��
&�����������}�qӂ'��p3�0�ӊRþ�~,���oSH�V&��\A(����z��帤���H�����ЊZr1���O��5���U��Q4{�pv~A�>'�����ܿm�tѱRVu�f��$I�R��p#΃��dy7�s�`bv�iBv�����p�T1���7��0`Θ0�QРs�BW���m��$��N�l���92!$��n���Ɲ�QQ�l?xn�0�����ڞ��*���z�*4lx%h8�D.�vr1��
Xu�`���6��n��� ��G۾:x�[�� =������[F�w���E�[ۤ�jl\��٬!l�zj`�%Clw	��
������o�t6�~K[��}��B۶�P U�hr��=F�n��vT�����!��D4+��%e�Q.sR�z�bċ�?!�B%+%%nz0��oiM��?+��ե�>[Hv �6b�
���v]T�4f��+ORP��2m���U<�e&.W�r�>��JT�i�<�s���S�`�,�B:�!ve�D�=/�P��a]ڰ�ł�}�_"�ր��3W-�����N��|]�#?�F���x嶎Ojs��M�O���2�Xn%j���с�=L�k��W��)֘�)ݜT!U���4|��.bf�mY�d�0%�WU!D��`�V=5��=�Tc�y��Ѩų��I~��Ms�g?N����AW���<��b�zB��AR>��ن]ku�]2)#�W�&�7�L�9��.t��ܠI_�A����!Af�L�@d����FjH���IJ�oeM2Mq�Rz�����v=��Ⱦ�h��Z����c5�X���������#6;K�?��l�k�������� �dxv1�m������7kd3���V|C��h��2�Y�������TQ����;��a��#o�s�L[p4�&�l�q>�-��p6�X�6���G�N-�	��L�!k��yp�l���hs������V�^uA�7��i1߃���<
��0���X��MS��9�5����}��~�7�E��͹=�>�dvAM�(��R:�'Q��M]t�@��'�#���9�'��>jFA�&�2�]�D|	3�*^��/�X�u���q]^�F��k�ш�cR�<��l%»�:�G.��#�qq3L��>cD'�H�0���5�<�T���"�O&wa�m��%h;FWv�Tv��.ք��H	�������W6��a!8*@�x�6�J���r��U<�a��.�Lb����O���kϝ���[X�V��l�2$����g�#��T�=D��rܥ{��/
�B�*����F�nrQ��U��JǅyX��`є�I���c"�(�� �#?�m!�Q�'��P0���>�=��1�x0jX�������T/���N�g���Am}'MӜD$R��">a�~TW�4?��TOu9�k�^5[��Z���@��1��%h���GW�*���HL֚��N���>Կ-���@��(�˨y�����s,3J����z�=G��^c 6\VR��_�e'ɗh��T�0��w�<+|��SL_��7�(�ɵT�l�֫3�\������@qqH	l+q�-�����8��R�#��]ut�!mbO��J����1$�7i��r�#��'