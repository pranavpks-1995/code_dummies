���RÝ�[�[�U.҉Q�%��(Ǯ�_8����~�����Y�z!&xS�.*���6���3f����A-��JN���������@�u��iP5n:MPն��&j�)�
��Sn�:J?��l?X�sz��\Egv}�UQD#�� 5�9�Y	j'�5i��|�o^��V>��t��c�%�$�� v���u��M�7`��l~5�-QSvm0�	�dƙ"͉�+���`[��7�ɸ��|ř�qK� ��/X����)%g�HK���p+�>��EՈ[;f�t��1R�ZY�FHH�� *�&�k����Q��r[׽���D.9�+v֤$�)Py8u��k�%9��D=�h�N[�e�C.�.�.K��3���̆ׯF]{Z�tTLڶ���nv�Rb�?'Qզ�2����<;G���	�Ȏשj�����k~��֟��=�3�,i�q�O��$�l[�^4��B�_������\�1��\a��ӷu�$Tzfh�0�w�CxB}������ib�i�W:z;���0�9Em��*)&Ǒ�����2�c㗇�ҬX��"dѯ����&����C��4�yz�r�����{39f�[�<[3wd�W*e#��M��<�Y<�)�'Ԟ
�:���#�Y��<�B�q�~������D�Gꔫ�Kfs~��Xl�����3W]C�px\l�!<>�.����aK4	9��!�P]!��Ov���(������wC�1}�U�j��
�5��[%���W|b���kC�)��@�>��	{_*���r�0��&�zϕ1�G2f�.W��=Xbԕ�&�:��#����=�g��ܹ�<�m����D�����g#p�%o��(X�/�^��h�'w������逋��(R����aG�ģ�kU�@ ����$PbW�Vj���n��to����e����u���p�)
�g��M9��~ut�'�C�k	�n�AEy����T3�b�v�A�7H���'_mhE�� �w!�H9ȶ6?���󾷍�)�$l'��,��p�5�="׉æ��w�:�Z�A�2zI�L|�^�)c��+ �B��_���mU������D�Nq��oY�������	��g*��1����l��?3qj�x��.K|QĊ%�S�Rnق��[�� b�N�ٯ*�k�X �zQ�܂��eO�Z�h˯�y5�[7g���+�A��U" 5���!2e����}�'u91vEvw9`��a�T��x g<�[]!P��m�L5~~�g�˾#�^�G�.�4$�� ��A�����Jk�����<��a`�%�Ɖ$ ,����
�t6��Paյ�w�q���Wbc��ъ�Q*��vҦY�p8�:�\�$i�L{�AQ�b�A�\�u+�ֻI,��P{�UI��G��*tO�-%9U�P�	��8���brz�OO��_;v)]�Ď�����<:����@�m�k7F�ya�Ja?:�̶�hy�Fpi���&�,�3'�*���!�FȞ`�%�H�9CI��Y�P��6T���yi�w.��}��F�{0ݬ�AaŐ��
4SU�=q
a�H��t��|��.�y�����9���;8�;����hi�r��b(�H��� �
��(c�����?&a�M��ʚ��	�*�P6`|�ꠁW�L	���-Z���J�Z0��?�9p�PУo j!��$:�aف�*��Y�ZG5;���X��\��^��Gɇ��:]��d����@R�)acWQ�<:Lȱ)*�:D��NX�ęV�w���~{L���)��e��@yKaZ�橀��eR�$�*Oj�[�]��c�p����X�{���\�l���zhYR���-��W�\�R�Ъ��m��(��Ig�]�G#�.�ja�&��P�U�z�)�n���0r$���Q��͓��(�UN��)�q���� I���_�F"z��4�]-���'�`�瘙�d$2?"g�Bǐ5~m��������S`��W��B>1
�Q���T��OLTЍQ�c�_��J��d?�����H N��=cg&H�1����ZXr��]r ���Q9-��[�/�C(kHJ�7D�LZ��U��K��y�/� �h<,�W^�I3���r�k��Y[Hk~�ZF#�d bV�����f4���LFb����3y-��F�*��:��ٴօ9�+�R�>s�q��#O;�[�Њ���u�S&�HH���$Q�CȊl|Ho�Kg���e+>y���6����O��H���}�N�R��>́�PuIm�s�Q!"!d�'�Nۈ�h?���k�S�����Hύ��I��0�¯��O�U���a�a
�[+{���ȉa��x[���U�ݓ��W�q=��q-k�}��,���L<��?���Ŧڎ:�D�G%Ǝ1C��(w|31?�(�+��M���UX�&�����&,��g�Y�rS����y�:�[X�F6���>�;
-a�Ԛ����p�XI�!XP&���ȅ����>�Q:�{��l�A��w���"��`�t8o�C���	Et_I�8�%qMIW!��7�c�	[�+���Pv
l[К/v�f^?J����B9Ӯ�D����ʋ���K�.4{��{���!�]�)����Jp��
]ą���`���@/��1�T�︂�����H�4���D��à]��>W�k�>�6gM6d�3�w	5E��;�/)���F���K�F�+i܆�FL/�;�I.���ur��	�+{��=�^�����9���������i��b�!@��)h%d\_��Ѫ��4�����	baq �W����X�� ?TA��r��2�^���Da2�)���1B(��t�qk�ᴱ(R��?6���t~���_�M��rrt�e�f(�M�ϊ�	����ψyc�#���!t� �^�v���n���X���)�嵰�g)�b�)��H�C�6>n�V�5k�'
"�O���q���Y����h�{Q��Sx�L|�r�g�y��>&(e��&v�%��<�2}uV�QzG�&7EW��oz
*J?F9��I�%0f[����6�e�4����VU�����(�@������'�K2�}8�7��U�>Fư�|��{�1݅�+e�Tu502>�� �T�Y\ř*�ꉍz"���ƒ$�����7�Qo���s�;Ll?��{��Q��Hs��+a��z>���4�V���1xS�V`�t�,����l��Q �Ro��k�1gdȍ }�4����_�"m_9��(��o��i���#�K!�ݤJ���K��x��O䝕����x���)N�rf��*;e2nG�p���Xlr�Ĝfyf���9��^�g��/ϔ���%�O�>�b�^@V�f��Cp��>2�Sr5y�9Ձ�FO^"U�g�b!��W�����u���]k�GGI��4^tH	���_���C�����݄�хK"+Ԟtz���Y�6�Ɩb7�<�^��4��Ƀ�]l�y���z�0N9+����|�A�&"�)��4æ��	Y!�����jR��(?a��?A
���^�E�%��rJ`�F����������'�-�s��5Qq�P@T�f��MY���\�5ݠ�W-�׸���Z��A�Ϙ�y��1d���}Vh�� ��$F�E�oA���0k���u� '��/�0���;A�y��I
_��
��QZ������U���r�Uρo�0���᠄Eh��[�F\�x�����+�g�}y1��;]}��W�0�];jn;X�@�m@�j9�x �΁si�@�H���[�L|�AT���˨���H�D�b� ���1Z�0�1W�D	!�/G4��Cc�[b��*�3�F�\iZm� 7��y�� Kl�O�#'�(ջ�J	B,��V֏�Wԭ�[D!�N� �J��h����ő�m穉P���-\��:}�4O�P\��V�ϒ]i>��a9�=��v��S5(�/9�L%�mq��5�������q�BNo{ 4,�1�(N�M?�&q]�,�ޘ=�T&��~�^$u��?��R{�9��$1�$�X�_@��=C�"��I�+v���#
���)��Ub_t����i�x�ye
���o��e�9����ߨ��������ʇ�PSb��>���Ӈ���{������麢�����T���,b׃���F���6d��WX�z�BOI��k�	�W:�f����b��Ea%�l>�)����]q[���$Q�ɾ���]z�:DLS�f��m�܇Wa�]�Lc����
�jSQ ���'��bMَ���P�E0����O������3���;��:Z2�4��h� r%�Nmw/X��O�{Ļ&s�'~��(p�"��܉~���.$��B�G8��˯�Ig���E��S�~՗�	��-'q���-���)��pT��N��tHmzXV9���k�0cS�[[1��KĀ��`�"<Ƽ%��i<�m���lռ%Bo��xh�N���ݤ��J@�&��Ԓ!z���F�t�ɋ*E�h���k~3 ��A+y�n/�vVbA���@˽*)'c��?���ǽ�B����
7� ��}\�u>3G�5ΰ�1IyTO��(��'�jX��4&<���8�� �LSv����/�I����{ �3��R���m��/��� ��%[_`\��G�ێؕ�R�z�"��F�a�?��Dpۉ6Wezl��'��{���sV�j�^ G����0Q,��O�ֺIo���b��PZ�r����ȎQ�p�eR#��$�T��K�'�qά��S)1)]�}��(OP|�ń��1��[>H"7o1PX�Ϻ��D�7�4y��?���G�6d��f��6�3�����Vt�N��%%�չ��!�(n��G�t�Y�N~qq�>rث&�Y��h�&�1�):����M���+����+�"棓-fm�֓�v���B}�����1���B*�r�vT�;^��h	��'�z{1{\�Ab���E�����v����3������G,h�˻����ZB*�qD�;������Q�-�,ԁ�4�=��N�T���D���u���3a�
٫�2;h4�dHu�J5�ଢ଼L}x/��i7F�5!�^$T޸���$���s�e�s��tja�)�Ǻ���D��>�,\6��?�=2wNe�ĕ�����Z��'�°���� aÇW�B`{�����w�;���D,�N��|]^�ƭ&몾�G�<��P۷N?��Ʃ���*�W�q;F���w9�Z;Ɨ�	�-�!�y�ͯ;�_�Lz.�wj�7���I؋*)���!��WR.fч4B�� ʛ����T��~�
��pt�������z=BbPTJ�10�ﳪ�b�)���ї�_T�d�h��̤�@{�������t�%@{T�c{��U�@k�� .H-�rO�"� q�
��Y�yW�G��MV�h)��M2"#k�B8Xכ�~��Ǖ[(�K}ʐ�.7�a˒~�w�����/���\��qoV��| (��c��U��t��j%�'K=ҿ�;����(�]L7S��J��x�zN�թZ�#fځ��n t��g���Jt���pWH�\У}��b�9R1(I|]��-u���Ň@��M��=s�)=�j$ = f���^j�k�^���1��Q�����v��u�w��
�Wlɲ�M��tф�d��*a�H�C��ʧ�Hj܊���m��cų'�@�,p7gy=�1�Ï�6<P]ϼ�#I�!J�I�Ά�s�?.\��3����"��~�l�d!�Ҝ���K�T�V�e�#��
�e�)���^7P�_�V?)͵]Ybá �``i�bm��)�h]L�G8��t�Qw`�/�y�B�9Ϥ~7���;���"`U��7�9������b�u��}&'����z�1����5,mC|T*=1%�����kU�cP�.1����F8#�������r����+,X�&��c�S�賋��p,�D˲�q�O
V�dQ�(P�',�ѻ�o4��Ca�lN����&��=������o�ڿ�s��2��6�h���V+{��a��l���tj��>��C��*���\��Ze�V��S9�FFM��^�i�����ˁ.J�#��E��6h����Jn��R�����Cu���]��Ԓ`@�2R��h�O��#�2��w<��:�hU@{�<Y(�!)/(O�t[M�v��׌D�Y�^�'V�91~���������5\:��fc-�s�i2��^Ō����T��Hƚ�+����bǠ���A�n�4���W�.v�L����o�pG]��I2f."���ѶG��;��]�@��rz���P��,��@���6>
�̷>�+�����9�/ߑd>����V6Xg��7���:��o��NBV,����aϝk�o��_3P�g��ҧ�|2������e×���;�)��x�w�3�.��c�[D8>��SCLW�)�pa�}�E���X�X\�� �w��7���C{z^��VK�#�h͂=2�W�$�I��U�v��:��V����5%�9�%j��b�?������/q+|P�OT��w�O	����EY�iYʰ-�uk��`��+�nx��Y�|�0�z���G�S���φh�������Kԍ��l̻i&Jj n*MOC��]aY�[��<B�7�cܡB���(��݆QQ��% �/r �h�/�� � LR!!�%Qո��.�����kR�q<�ҽK�j��걯yH�]�ǔ�c�)<3�X�"2�X�q��� ,Wmb��pt�RΐC��;�F�=�8,אO�)�!��b̸��ީ�s��쫞.�_��1��C&��hq�	p�R����s����W���L�e?9ͤn�:b]c^U�ys"bzqj��Mv���!΀X�%�;�� ���a���TFl7�h@�K�i�B
΃|)�
����|�s��'y��Ҿ���ew��5o;�I�ś�Zn�~���]�~*���q3��J�<����9c��k!E]&��@d�}�@�iUhI���&2��*����F�*b�} ����xA���?����0Λc�v�������m��
s�x:M��zV��	��~�HK���J�S�\�F���@q$!o���3I�|����̘� �D��
�'xh�[Zt(�Q�0����y���ӟNp�Zƽ~(���~-H�ژ�����̙ڋ(��={5N���}b��gwy�[0 R�c����7Њ*q�\�3e ��֕�� �+iU(�X�xg̜R'��a1��r\���D^��dI����h+��s�g�y� �*�A��7���onޢ]ڧ?�#ĩ�)��m�C&A���������i?�h��Չ�=��c/�C��E�XԼ~"�%��Y�1S��;�Ț��82�*�_�ܞ���ȍ��FNy.!`5+2�+�ᑓ�H3S�I�5����8.\�ūc�9������j��5�~�V��	�؏�h�bS���1��6��ZhmU֤�5�̨����=B��O�"�
������-�v~=��P���۵��.������t{ɨ�&���JHe����E��/����eܬ{w��P2|�������J�%-Wh��6D��e����GY��Nk5�J�%򆓗}��W�`��
h�6W4V��k+�%|�{{	��5){.V�����+��c�?��ũ��<�KO����������&Ώ��ފ���7�%���xQ�r��.�/����'�h��?,������-�
��$_��LN�ce�f�Ǖ-E4]�&Y���upWKt�V��J͇0����T�M/�b�����Ҟ��l�t	)�^xV~�Q�:5�s��!��+L#��/׻nő���Ըz�9���:�hד��
���(�|5(����qBU�6�a�U���v�)Q����7^���MS�ejcw��̒J��;Yu����wg���ELy��ET�b���k-o��~�
`��R)��N��-=�|����b3�D�Iȯ�����fQ������M�(\�* ����n���K�;�?�����'I1�-p�{mH�H��`{!Ҩ�	�<�A�1@p�K0�L%~R��sgl���_�K���`!/�u���Ǘ�~����9BPW�	/%�Z�9�}����fuQ�U�P��I��}5�KZ��|//���C�.q�x�oh�����4�  	�R��'fJ 3���Pΐ�L�j�l/������I�l'|+��,4y����-���$'���w|κ���6��!�X�����WD·B����.�sD6��j"���6V4�TF����vǧY̷YK�Z�A��2����ם�����1zHکĆ!�SH�V��Tow�2֯u��jGm�Q�/rU�]�J��yCh8���|�}�`G���`HJ�@��ev�9��w(�,�J��+'�����>!s�C"m�d|�u%��J�j�}F�H}[�;|l ]`F,Dqh�q,�+�VfHI�s���QT��᥁��)�@�3�i?���B��r¼|b�@g���R>[YpgT��ag�*�n|���9U�α�ʱ�^(Z�8�(Gu�X�����.��B�Y�Pl��z�����P��eoj{�6o%�Z��J(	<���uR�Vw�k�yEz��V?���v �Ĳ��8������e��\��)%�	;�H��]6 ���U����f��g+Oy��6��N:`�}i�c�����7uODAz��I軺 ����`^� ��I�ir��g��`<�n_Dy��	�y�GO�l�Uw��D��G:LN��+PRvF��
�����0�P�r�h`��4-}�t� Ӝ=�4޾��x�J���h�9~�!�#i
���BV��Wɖ���U;��7n�b�8�W��m�2��J�/�٘9��`�w��AS�}���Fh�w^�����c���{Y����H
!�����J��Z�9��&L�u[b�[�(t�v���X��%�u���H�G�*�Y<��?5k����r~N�d�}�b�{�,��+!�2j��p�������5�%(��64�Hڱw�T I �=rZ�o$�^��������k�l[�B��;27�B�N�e�9<1É&�O�� �c��s"4�g��A�3S�`_'?,�����ǉ�g<��� �6��,3�YD}n��c����%�5fd�S����	}��w����
ʪ�{�d	�QR��.Ԫ'A���������ɏ˾�5�'�+�#n���73C�?��$yd����͎N6��ڦ�;8�vH�&�6 ���o��,� �%�M���ʽ��{x��"L�><�V��9!3��P1a��8�/|)Y�L����w]h7rפW�X�L<#�FqM�^OI�o�[p>f����C���S�D����Rj�Bx:"�βC$$�M�:������'M�gnk���"}q����	���Ve�<71>clx�Y�z��#J�����`�n=d��W����Rʂ���砞�2{"���O����.���ǿ�����?+�c��{��n)�H	�����F4&��ҭ�]U�q��.�'��V��|��S9�Գ�㚱Y^�P�L��/ޤ����8��D��&iu��[��8)�bZLl�1�q3�)��nM���صA^I glM���V�w������� �����t{����Hd� W ���?=x:�F����s�_�B��u�3R8#�G�}s�>i #r���L�|<�X���}pp��y��Ak������Y3��0�oF�K��U�R� ��́�4�b��l`���v�i>��U�Gh;ئʩ9��`�ňk)u���1��eN V��׈=�� {|��L�E(e+ͅ]�&�a��}����i�i{1i�{�1+HԽ�;(#me�Y�����#��|^�G��`Ç�#�,5�5�':�	��'����&a^8̃x�;�t���?�ҵX轼�
��z�@=Ec4�M����-�Yx�s�z9�)s;D��02dl���mp���i	�Dh��>nFr�=�R����"DnڬU�(�5�8��h%�ˍX���ˀ�3��5�EI=�`*L�.ç丧3o�J��&���:��x����7���Ipl���|�F�ә�6��dP{O\6���o���^؂����GZ�@��A�71����>�m�`��*hǨ��>�ȉ�/ַ�asN+����9������p�� �g�6�w���	�Am���86BI�ᣥ���$s���CVM�8xE쪇~ڊ(>��ޅB�$!����tæ���F�C�+���^��c���{rP��Q�wh��n/H�fd\����F�r,q9?�^�ʴ�G&�WҌ�_t��}v����S�$iF=&o���;J��ۼg|��#�f�č��!�<÷�5�����	�{�4�?TE	��b[2�!���ӫe�W#{]��9�;��)$�t�k�T�b��ꨂA�^)!ȜJ�]*�>B=K&Ⱦ��.��hUB*����������=�BGż!U�aV`4�P(�cI6�u�kxC�A�s��&X�ĉ����rm3-r�)���h�����+�ѭ�+�8(�vEٛ���/N�|��x?~�,�E 3��� �Z3lw��x/X.����b۪/^�؆�2Ҫ�Bg���:�Nþ�	�.P��Å�
>
�iR?�m�N"6t��'܆$�D���w�QҤcr[j���J� .'�ݦ�K}^�!��!R��P���4���V�gc�ܥ�V���JʟP�=�7�Mr.>\=�NkH�n3h�|����fgp��9#����Lzj3��#� *7s�ç����k£�m�η���\e#0�1{�ׇj����[蛀IG�Ӷ(󬄎��6����=jpu�l�R��pHv�逶�Ea�z/Lӭ����~�ކ���Z�h�@�u�MUI�Q�A�����	��^�Ӟ(��Ht zrW_�H����R[wq9c�#����w�&��T+���T�;�Hdd�:޺SĦ�r��}w�.���k���h6/K�������!p�
��/����x��-�7�  ���W�GWVQN��6潯9���?�a���H�X��W�U�>�Y��ߝ���p����-�j\�h�'�N��7���s�E%�؄��h����\�l0g%Y��f$k9��［"6��c�̙�����-�E�f1�� Mѧ�l�j�����0L�?��V[��MN�b���痼/g��s��ow�Y�n�ӫ�G�#H2�A.�����	Ο�{��}��Ԁ�z��c�)-dCI�l	��'#L�e���fz�/!���=�J�û�7$�D��6/��w?�Y�;�P�L�hɼ���ӌ�qķP�0�k���u�qF�[�r����&���*e�'z�~�6Bg�VEaS�����h� �
�X��fr�X�i�L�	X��C���F�3-�
Xa+ބr���ʘu�#�����_H��ț��4Z�G���po< �T����mq��|Y���l|ص*�>�����A3VҶ˰����:]K���?��9�;A���G��0S��c�w�q�F=�%Ϛ�X���}Me��ãv��$����u�;�����J�tf�
"�P�n2��F����u�'�r�����[z"nu��&KB� �?e�.wVʊ� 5(C�J�� E��E���{�<����\���b-���	��m�����8��;��A�2R�q�)��s�;����1��H�/˖�?�
�b��c)��Y�(�P�MBE�Ұ����oE��T��gu\��6����J8������d�m�֮�w����`1�a�E��ؑɽ*9����n\A�f��9
qs��S"��U��S��4��6{{�2������M��ȣ*�aI'.uUZ4c�fOt���k��r��_X��Q�nw.I0���6����*��UU�+Fet僴d�\�^�.��W��3�dikK���A������7}(^�;˨E ��d�Jː�q���*Hch������i� �챊�pT���L��j+�-��
��xT6���u|s@h��D�n��_#`�@�i��c��lT��g%���#Z�(/yW��ǐ=a�+�2�.*�5�9��f�i�z'HO1� �~��=|&�V�!�DSk�>>��1��n#�.L�#36�0-/g�4��b�bT�{ʎ�԰c����V��(�W��Ί"s�R>+��$�_k����Kd}��\?.,*f�:1��=� <��!U�_kSR��W��+�c}<����ܟ��+�顐�Jw�2���B���@��=~�*,d����S+���U�}>-���9�����v���M�;��n�A �Qö$$]�n��![>|)���2)
%Hm|�(�{A�vn�TyB��޹K�zUO=|�EY+�k����UC����~t��A@�s_�p�1d{H�.�Z�P*�	���
����B~�ä,�L"�����;�by���