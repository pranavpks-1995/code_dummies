�>C���2\M�����.���Î{A��@v%�t�^�r&��B4����P��_n�z�>%c��B')0��nr�
Mk�u�a8��CY�H  Q�'U_q��z�~f��pd`S��͂���"?�/�r ���8�̊��Z��0�9��ӷ3��n0$�q��+���^�pS�6@�ٖ{�_Ċ�DZ������8-LLB�㚣e�c��V���HpĔ��5���������/�̀/��_5�Р[�F�B*��)=]�-[Y�7Ar�Y�˸Z�
��~8gNd�3:)�8#5^�i��;��ٝ ����P�w*��d�_��o���5k�d��;dܷs8���q������c�C��:��P�>�g9�rf�띢��7�(l+�8�'_�x������`��Ü7o�!C�/J��?�(�v~њ����� �b�Ӭ�}�Zn��y0�k3J�n����Ju��i��m�4��p������Y}��9��)Է�ml��$����h� �É�j����\���-�a�L�-�8�0��T��1l�k���1z������yi ��D��{}Ru����	>ৃo����n�B���Lߪ|0���uj�J9����]煊÷O��_�5������LD454�閇C��dt��Ud_0|n:n��5@����L	A����i(1v��VS�*0%�ׅb�����W�:u]R9 c�in1�y��7m�V�u�w��[��y�Z�+�̸*�~��՛��DEj�㓲�٘l��8{W(с�<��\�VQ��h..�(A�.��O��X���iS'@0��އ'W|rG�p]E��Q�����>I��[ �GƵ��3?�3�CC`6�������DoF��D�ɢ�՞���M��4���7� o����4��VV3�������5��RA#�t)w����B<��  4 �f�U}"�F5F���:$��u|��k�Q���lk��w�GD�nKA�$��f3�>�&*�]��M��K���NN���� u ��[�f�oY8������긽���
J�o�J�k���<2��O�I�L�0�g��2ǧ��m��`��N���g�4��z�b<iB�I�+�t�O`G�MyQX�����PM#�Oi|]`�X/l���,W.Kľ/k���H2P<6�y�m��#��j�s5��׷<�H�+�z�̠��pq'ڝk|7�6eM���녪U�- �k�`˥�HV��,u��uFƗȵꕉr%C�[w�Sߟ1ui�%��7i�Y�֮���3 �����k��Kz@�V�Ծ#+oͭ�8|QO�^�x�mZ��T*�(��0Tɰqh�`��!��m]m��%`����	}L੝�@��H��!(�*����縵m��Lˑ�V�n�h�M�K��
�$��z4EPUV�[B}-��M��(˧yY���jk[<��V�]܄���o#9��E���|�t?:)���˽f~�Y�M�d�r�:4$����Y��B-�   % �ԝ}"�F�� ю�ڢ�6*/~R���g�L�+��
��t�Z�^����$S�����9�������B�����M=�D��`��jv�!���������6!��.�j�x��e��׋����Csn3�}�.��PLɬ���[�y���*cN�������@��"۱��s$�m2��K,��%~4k#�,��Lt�9Ә^_S�5v�3�>~ڌ�ʁ�ω�")Rߕ��u��yV�ã�����c1-�$|�쓄��z�|ocA��]R��qg�IR�.4�.y
U�6�e=*Ь��몟��Br�����U��v��<ΰU2L�o��M�V�-�v�\T�2z`��aKh��r���U��;6'М�?W�&��R�,��-�8 XR�D��������p��z���l/��ݓ-�T��]G�(@���{<�F�ׯw�!h��\F^�{M���
�����0[���?_���y�G�P&�*��� K�게��R�����f&@�s+*%G<j�Ɩ1FÙ$�N��y~�Aϟ���Z@.�tN������AS�r   K ��-���:0�$�
�®$���p,S�]0��M�e�@����xgl3s��v=�X�g=�6&�>�Eҩ�H B���|2���yZx�RA�6(��an�	�i"�mam.�z��*�<���.?�BƋKSKw�V-=�����2�k��y�D&����ɍ�H;?&�Ez�8��p���鶺�βJ޹X�S��Y��.�_��]�U���
LWP��Z�fN<q�a������zs���p�i������'_���s
 @_��nG(�W2���U�<"��@ޞ�D�JB���F#�A3�f`)S`�'�|U���J����g$x�v�ș�(�����, ...that collects orchids
or has a lot of birds.���Ew�f��������!�����@("��� !)�Y*���eʼ��J7>S"�ԊE3�B��1���x[�K��X��ki�
[��rX��Dv�
�09y�k{�_��H��6�%����3aM�,��V�&tp�&�ο)��嘡�E� �"I(>B��f���=-���  !����*P�p� XtY�kQ�  �A& <B��|��r���{9���f���!i#�3��S".�͟m�[U���+�v����V4n�H蟽جJ+ҿ�T\A>��k	Ӣ�`Qs �!y�p�)�-G� �A=f�~x��B�����
y�  !��aHAN�QF�H�l���s����8��'H���јH���9Ʌ�r�(��,��W��-e�( ���(��=}��{ ��*Q��b�1eT�������{�;�竀T��yA����d� ��l��6�f����N3p��  !��`F�a@�"Ex� ��I��x���}";�'z�0b�_Tv[�H&���h�-�Q�b�.��rxΔ���Lձ�n~e���ʿ΋-���D4ڴ��k�7�P
w7
���0�wl��(���������4UM=��H�R)n��r5��a���&M!��p�uM��U�US"Ĥ��>R� `   ` !�
HX�a@D.)u   ������Q]�MҕL^%��&���	�4�o��֛+\�WZ�d��	'/���/�L��b�!��~��6uMu��?
�o:ޱ�ED���6�^����ҿ�Nt����^l3:m�&X|}l ���Ӥ
_�Wk��J/��     �!���'" �B��vn��*۩���d�pk��g`T������_���A�?���~�4�V���"�������P�N��$���}% �9�bǐ�q�*#��wpu�h�ύrQS?���S[ٳ���e*	� ۂy�}.�K��^b 4���S���ʉ��2���0    p!��**A@  	@����'ºEδ�Y��0�e�V6  �U��kVڭTN</�z��0OM��1(��
r�Ϥ���G\a�ԿY%�I�2@�eY�&q]�_{�^|� %`h��$ X ��8���	ᑗj��B4� 8�m+���w?�ߎ�>�OL)�~�1����Fn����IX��     !)��	���P�V(2myE;j�(��n�E�7��g�K0BH�ͨ'�$0��c�p�S)�ֿ|��P�T{�FY�)���qv����CT��8���Ej��K2���T�S_�Ro��A���O�Fȹ1{Ԯq���b;Eb���b�@�@  ��ŷ�[��٣]�9w�H   HB^�% R�4��S�u'qԇ�     8�O{�l   sԠ�����c���y�Gr�N�8�9�4hT�4B��̆�a8Qo$,�Q?���kj��7��b2����D��6u��M8���3ixA��gz���C���p&c��fmBP�H�X��M�0�C	WUU2ϨT�N�QP-- ���Ǫ�$�F8�:-��@b���P�ي!�;��-�,<�*k�����p �f������]�V��S���e}Ñ�^�33����r\Y%(�`�sa�����Ns~�qB�!��������ʹ3����<�T�z�j���{�nh�G�4a���$a��Pa]7��P��5����u8���^��<
�o0��,p���X$��%4�b��-�S��/�K(?��F�	ݓ	Y��V��]x���?���̿�x�^�p���(];�\q�V����kOc���ۆ����l�ox䶹��Mb.w����b�eYH�6v��|��"Oó����q�6j:FX��LX�e�~v���@#Y ;���;�?��/�u��ޯ��+3|\���+������[�u{`<�G��ĹL4s��ZJ�x��l
�c��L���(�%�D��c�l����h���?�d��5���!��ʎ�LpD��+p�E��E��ͱ'`Dxi�9���B��2�P��G�G�o����	"���8Vg%��N�2����V�<�y��r~&�������"�7�N`�J�X`����<�W�Ͳu5�Y��ؑ���A�#�m��d��T��y�_g��ˍ-``ez2�����B�ʳ�Y36E�}�0'��]NOl��h�e�㘕Ir�H�����JS�����pF縎 ��� {m`�=����Sɱ_��#�_����
"X^:/*H%�kx[8�cݟ�5���}k��j�Ǎ�k���"��!����^SkrQ������Qrщ@L�{?;Q�JHz"�!}!D��_� �?,� �������mN;�J����{�1�l�*/y�h����=�vf/�@�l0}�ƶ(.@�q/E����l���`BOϻ��¬g�!'D��h
��� x�{�'M�����P�Lq��5)0��6��ָp:И�ǙV���-�Ǝ��9��%\�N���ꝍ�]�tK�!ƨ>ӝk�ę0D�� O�.���?L���.������q�p�Μ����+`LΗu�;,�������˅D��&�1O�B�C���{U+�������4�fd�	p�m�k�LN�N�r�oK���c�d�=��@n�����ձ?��"�>��"��$|֏HZ��|�+]��d�>M�~��̬���y$��тޏ�QZ�K�^J�I��RKLX0�'\������q�s�+)��*Za�pi+��@<��]cG+X9��W�r!�xф!�\ɰ�?"�w���r���Q�k�� D2Ǭ�Y �@g��|U@x���K��g�YY,i"Si��j��U�� �7Ɔ!Qv:��U+��E:��u��"�� �䨜��ߑ=�I�T��^]����	+d�.OrA��#��!��fpe��� v$C=v`ܑ��6�_���q�m��a����Qd�НxP]<�O�;:{��d�Cs
���(j�x	3��H����H�&_�8ĖQ�A��s�$����y���gJ�أ�Y�@in��=Zm\ߢ���`�i�����RX�2HG�{�l�ڠ��Z�#)�!�s�h}\"�9��ޡӯ�`�t�}	��~�0}����G�
�'dx�A�$ܓ-iۙKz�[ޘ֮�<*LR�ee�T�Wl7d6~��ˑ F��o��Uv�s#c�<ĵu�*W���Ƒ��I'E\���ثQ�^ڼυ*�?�ѿ��r�M?��9C6X0l�Є�Ϗj+2�C�íey�&��$���:C�uޗ��Miq5q���Bo�k���
h��g�f䋥f�gZ/�9_-ߩ�h 4xxP�3Kb$ܤ�H
d������/J����&�H _	Zz�����.��Οi\<�Kx+8�;���ݝNT��*V���ۍ�}�$���HA�o">���eJT}c��Z��L�m ��?�G�A��;����)XC9�Z�<�F)�4o��{�����.���+��C�������{�� ~1�~��fi$Ѧ�Z�h�@(+J���T@�Z0��-7�hy��]-Y3kTm��[\�z�x�XQw�}7n�/��%��&u�:k�*���{xr�� �ə��cAt��?�{�*�.wp�;NR+i`4"K�:������_SUh�%)�A��̦�J�'��k6�w�AY�8(���ޙ��9{�U�Q�h���c��Zo;�����0l+`sY���=��&k�Nz��=�����A �\�j%�����i�Obcr�֔�b	-���`��n���{#��A�� ���^|D��h��N��6�n~[��a�NSk��@�I6�6���̮���|qe/�w|�c�|F�u�7'1N���!��3�$Ny���5��ħ��R�H��W��4�Ԋi�&�f$��ȕ�oD�!��|�[�e<�YE���(��)�����l�=�	�se��Ӡ�T�Չ�n��+WlI�����w��*e��s��h���h���%��;=i�er���M�8~.!��_�ѳ���A���������b>ӗē��i�6-�ؾ�¸�3x�
����3��5����p�����$�撃1�>R,s�*���!HB!�7���aG�y6�nB��L�ڢ5����ӂ#�_���w�JLM}~Y�3(�d��c�B�f�f]��M+!X�OL.��ȣɮ�S@�X�]�F؅�$w���
|���1¯��6L�N{�v��l��T���z4c�y;A
��И�2�H,�zJ��f&F��ɹ��n��ތ���j��ٞP,���,�nf��`,)�&UV:i3-�ʻk�7@�i�V�<��a���A��{ôQ��,vN>쑡�滒vfUw:u�#�
IA�VɎ%�y^F�@�?u35��O�q��ry%,�
�Gc$���Hz���	��AQ}� ����h+g�~�-x=%D��,O� ?E7�ӿF�.y#R�9��&�9�+9Dg�e�z� id�5��σ�����$���gH�s�ʓE����֘S�A�n�*�^����a��ve:���߉�.|R��嬘7﹆����<���g��&jS ��S=ʭO=Ь�P��J�ZA�F�Σ$�8�F��1�K*+FlGf����"���~� �(}>Az��-�щ�6���fty�����T���l�6S
iHv����Q���!���`��9�ӿ�]Sb=�Z�bb��xF��wך�Lچa���]J�'(�U�w"�ࣅ_��}"xN��`MA���\�՚�&�lqa	Z*�63��VV7�%��ky������<���^��MF��W�3��Tmwe9Ue$%hL���D*ؗ�o-��MK�1m��G�����2]ϫ��"%O�h�8B��n�0 �	�;ڇ�F�@}�p����V��p���e�]��k�}6� N���*2/Y�qK��5��x�	4ɓρ�RS򲅓����z�J�N����v�j�W�E���3c2D� ?X�2��)/Or��u���6��G
�R>*x�2��1g
Y����1\�0�]q(�y�dg_���xH�	���G��`6�T���0;҂@"��%�G�\���1��,f��b���C$�͕���������z��	�p�� �-��m��塑�@a<�)�H�)��B���`6��_^��\�N�V�{Pu&-~�D�83��݀.
5"U��ܫ%��1Sw8�\}Ċg�UE��|!W��7|��ii�k���d��%-p[8��ÖY!u�E��'Cr	k\�;��v�ܜ�������8��ԯ�
�0\��V�0�D��  ��B'W_q��R���{����;�H\�n'J�'��n2��ڴdAm�t��
�u�r;"E��F#�n��O8���\a^��:�}��c��hD����̝Z9���`o�Os��G�K�{��h�ڼ�KH�����y�PE������7�Hl�Jy:���b��a��~�t�����4�,���J�QRn���¹�5 _��$�3��&@�s�RvO�-��m�*WA�������(�`Vs�0�GX4�|�b�:���8�^�_���Dg�n�җ+����(��/̝g�����ފb���m��rUP����ݸ<����@�
�{��'�{���o�!Љ��J����yc�)���{�C�R�7F�����4!������T𹂠�f�9��l�n�w�R#�>/@�����"0��Q�#�C ��WϒԸM_`���t���?ߙiMe���u���J,���o���Y����X��SL�VMj5z=�\��Q�W�p\퓗�6��i�O�
�(�����N� ����6KMUa��H�HVm-��Y�=��	)���ms:R�t�3���l��(�U|d�\D�U�V��P���l=1�ה��k�Ԝ�I��8pE{)]�nU��]+�nZ���2���b�Q=Htx�1��t��!�}U�H�NJ���o� �ha�62��:�jzz���|�0����F$�;�*�M"lP8>�����u{��ī/�V�L����/��)�m�h��@�e���y-u݉<�w=}!C��3��"�	rF�l̓_)�{��0�>yE������
�3y�̅�R'��R�Xg�V�e���?*?�M����Av���0%�v;��o��H������q܇�,�)p�>��[�Zu4{���Ȓ��߷}V}�s��y�h�(��g��*-�"�a�)u�&J�Q�Э��_h��~qgA��A�����%�`����u%�M$9dj��5p��q;,Kq�����������;chD/r,������q�P���
�cۓ�h��O�D��$̲0�g��;��^ܡz���a�í���"ѻ�(� �Cx�jk6��1ð�ڱgH2-�\.��=��	��0%02�~��<>�L!
d��(���h-7k���b���xܚ��� [�[}�f��!5��?�(�����0��Jf��c|�,�A�+���B:��  2 ��U�s�Ϫ\�rfm@�Z�z�Y�3gi4N�	{���.�T&�Y4�C��6E�� ����8EڨԾ)
�K�?���7L�;�r{�HC���� �ˑ�p�rǲ�C�]|d%��ؘ��4�};#�Θ����op@!<��8���N���з1����8��\.�)O�~��c*�.]`ss�^�<���[_|6��v��/�6�P3$aQ�r��gS��Ճ@;�(�a������ׄ�0{�t�A�-�`Y��@�<9�w��#¦��T�dS��ى�T�f� ���q<��|-p�%��2��wE��}����, l*r#p�6�/��<���_��}^�9X�í�GNn�*�y��7��.-�og�a���5&��^~�����O��˙��) ,ԇK�*x;�����*����C�詭Re��y��E/����$���,���vd�vș���7�~O� �V<�ڮ��ke:�c��6>����P8%-
��D�Il���.B@��j��1C��}_�~�\L�c
h�e���֤E~�֙��3Ft�����:s��⪶�C>�9�B7��   / �&�u�t�L�t���,@r�B����-���8�t�d
��6ZӇA�F��@lX�8<�����*�H�Y�qoy:�˔�|2���`	�#���"�H���j�a.�z�4l򨠠=���k�ܡՊ��^�-�EYg�W��:Ȍ��:�����;;�|��1T+^���q�Dl���ck<IUc<���擕����G�a�SH/�u���� �,��!�P���X�a�F|Q
5m��<%F:�)4��Pج�~��'�ITIH1؉x-=�>��g�Q{G; ����Q�?��SISZ#&L��3Pa�����T�;�q�5���������`Ȭ"r'P"O�(��]~5Q���#V54:��s(�vEy�I@2�;� [#����6�<��6�lƦ�Xz�b�u�"E�|<U�ˏ��\e��X
V�I{�����/#u���-�w�n���i��D��⮿3���1rK��R(�k>�j����E�r�Ѡ�R~����8��#�����{)L�^@!e�U�K���5(���ɋQ�� ��])�㈣Bg�B   _ �b-���Ö^m߫8���[�'��KRMG<�%+ƟW!%D"��X�Pk��g�8yj�4{�J@:���
l����3���$4.� �_@ ��)�����|{�JAB�^C�Ze�y�͋% _�2)zg���N��3�ݿ�j�)^��~��:� k,�v3�yM>��5Ț�7�}���j�c�w��𹡖E���Uf�,U�(R�}�A3y�g�ro=���A�~*����!w>ne�$b=z3�&�qje���7�&ozZ�J����UN9����~�ʡ�k��o������T�wK4�yt�Ri���0���X0o�]�ׯ	�͈ݗ���MH���b	�U;��-֞�� ��0���\
��݃\��YαVkp��X����:Z�7O�g2��1�oB�\�4�dbi<��ۛ �X��2wuG�/�a������"��ʫ��6�έ?�"Sr&�o��*{h��j�͋w[��HR�"h3��ޗx����x�\&R��'�R~W�ńܳ�� �M[��ө�����b&5ў;�T�A�C��v�'k��Ι��dI�l�+W�=�,I�!_���i�+��b`��K���$�Nd�=   \�Ȳ���C�� �����}��g? ���m>xq��Hbk7"��vqy[=HF�|���>��тiGc%N/4�l��_95S%;a\�:����`��N�!� Yҝ7DR��p�ꦘ�̥3
��X��z���3�F�
fp��Ʈ���8��6.8��럘�ꈅu