����r1�:�*��R�I��h����8o���|E�L����%�튨MB壮[I5z�m�Z��:�s��~i�SӔК�6v�ο�����:̱�� j;<�
b����:"�'0|�}m�8��a@������mH�f��@��X�1c��h�+�@��Z��U"Ɇ?uЌ)Ɓ�{[&���r�(Sh�ng�+�P�?�z��Tx�>���<o���x���A���y}y�������4L�/N���v|��<���� Q�%\,7���m#�;:���:�����G��&�:��*�A�!y\6:<�|UͬukϚ�%�W�5�0��GژP��=	�V����ꏒ♻9 ��u�o������]K8�'�!�����0|�/iz	�03��2ȉ�Fu֭zËH��_����M�t���V��i���BtS������G-/U$��5�ޣ��8#�xEuΚ��7 �!�I��z0ٹ����\R�����pz����l�.�GZ(�j��O]zKe���4�}!�E��9�z��>dc8���Y�
~�h�����bJ��M��W�#t�b��D��o�(�2�vǲ�3V���gE򧷴)�g�3��Na�F�X��a��l3��V�W�A)��ح�"4�\8�����_h�ȶ;f�W]�3u�N�4
�:��Oe����&n��J�s�|�2':y����<��)�<��n�^~�z�Ch�Kk/9����ݬ��^��K�sd��>�QGі%�"]>Ň^�%�n�]�p���?�V6���*6<�)ta@&�Db!�h鬹3�˜�}�u��K��PI�#b�F���+��R?��q
@{�(��?5�Y[���_�Op��{���6�
��k�{}��^v�e�[:#n���
w�`����%�G}��_q�u��9����ͨ��4��-H��Lՙ�;�5��׽1 ����|�GĘ�0�G�c�s�(Ȇ���dra�PɆĎ_�FB'�D�-jo��[e�U�p)��*�&Y�I�JF�_�!�����]�;�S!Ս:e܉��xh��������|���W�ң@��Zb2���X��:�:ZYXz�F^W�vR.IT:�眛͊���Q>�	��2a���g�N5ր�������x�=	�� WJ6~�q��8��Pc#�"��hz��G'�r�͑��ݮ��0(�6������P7|.��W5�X:��\��-:�тYqR$��m�۴���:��u���������0�a��M� qM��˴*����(�I����I8 ��U�M���x�Z'��tU���l��#��ZnJF���4l��} j�K'k5��_~(�n��x]!�h��
r�x���)����)�(;%\��2�# ����=��f'#�|x:g�zW�1֧ZT�L����[�wR.c0�r�~��5K ��@m�������Y��N
��x���-��!?���q��]��L����BC��m��k���7^�S<G��tf;�
b�e
9 ��2;��p̐���+-F\�!|��K}2"���_~T�qQ�6b=�}Ð%�?DfD뇂����P�f�y�C g��@`�G�B#������`��o2�D4�Śâ�}
H5~�|C��,�R*�K�Fyq wz����G���kDW�{�#
�����Gx]��3}�Z��͔Fbu���2��$��5=����n������+S��:�Y��~ϒ�:ϱ���MxEL#�ީ/,�ET?K����2"d1��*���<^M�FG���B?!=�MD�\^U����4$jn���p`*-���rbLG��4�qș�\�S��ޫ���C�8�KWj�DK��Eԗ���7�����G��z�ݑFp]2<��
�]%��p��Wa�%�s�Jx��j��xO�͸0��J�ۤ�+I���Hͺ��� �q$&lQs���t{-�;�$v32��� �ʹ쎋@n �**}����x�(���ăx��BT�#yS�w�+�T�m���M)�ୟ��q��"�jI�"*��G��:��&���T�\�GC��N�{�1�DY��5�J��BPv8y�K�r�|Vn�՜߮��v~ Y3u�{�8هC�IȘ+!���{\�U(K!��<Ds�#1��ppU)��)�B	���S�\��t�Tm�ÃD���ye8T�ƥ����;�+���y��vL�*v8:K�j��[Z]M ��Mhs9�Yk=�^p1�8��%�('�b�%�,ލ�t���h1�H_I�,��Gbf��1=���H���T'�QB���5��4�t|s�'䧒���5�+���,������\���]�]J����V�o�z�sN\����7���Ht��f��퐖ދ�zNoDK�t3)����{�Xy�-��t�i�-�4�r�#K�-�k����6��~TQ�3�-k�Ei�3�4��2	���u��q,H�9�a��`�������;��������hBu���Q��/����Lm�� b�)/Q�b��[��P���ƛ%W� �ynNoi˫3�{C�b��3�v�̃h&�� �:"ȝ��=b.PNO��7��u�4�c�C"�n�ێ�V���Y�� Pˀ�;�xj�H	
���9X��a�L���p�za�f5\\�D�tzĚሩr ��q����U@n8C9-���`�IXhf��Su�W�z�;�D�Jv,��R4)D�X]����R V,X�+�#jh3��>!-�My!�Q-�m�����J9v=8��]ey�P���2���<�Ja���ŭ�_���ͬ�z4��&�?ض:Z�(�#�lyE�t�ⲉ*\�C4n���D|ѫU80��,�$A:uF6�F� �m�e���d�!e�[�k��#W��7�*�\�^����%�)�ig���T�H�JD;�0*�A܊pVULy��?�;�ʯ�%���= �:4�_���;0B^��|ۜ���r�t���F�=�7�<P�a�o�LƇ	���(�~C�8�?���kx�H��J���`�*o]5z�3A��bf���ʿ�$�֜��,���58��'��؞�"��d�l�����$�
����ܗw��	`��񪥝s����.�k���8XE`����G�^�L�|����2�EfWOcF̥瓭��ۻ�|Ծ7/B���zS�%����B�谓	/C�,5�R��^ߎΗɚKpa7�צ���X}��[��0��w��6շ{��[�����(F�1;��ZU���d�L�B����?Yn���誰�>�Z�����B�2͞�ezI�;r��1�,���_�Gs�d�dΌ����A�����bk�y�&��6.���b�Sb�{��j,�gd������=d�@�����Z"id&-uA?M5;�?�=��:0*D����K&�9�eC`n
��ITa��й;�m�7������@v� �Mݿv��T��A����ې�H���'q BY��~�|� WW!>��	�(�"]��(^��׶5 *���+�sw�2E.)mW�	�Z��v�e��Jҷ����ظ�����j�g�ԯ$�,^0iPJr��3Z��-A
P����]�i �]�0j����a�(���a%VIs��Qɻ=ÒmdS�J)�c��8H62�6,�	�=$[�u�q)/C#[��=#�G����O�5�rw�GFHbg��+x�SiϠ�����Wt4��b�,�*l�x�n��� }�bc��3L���x}��}6q$.d �{[�Xu͚e�Y� �p�J��r�r8/�Uũ�G�	�Y��g�����B@�������X[W�En\`n�C�����w�t��4�冐t
��j�?�-�&T�����$�]�0a)b�.KK���Q���]>H����ǁ����-�|��|�-���JB�Zܤ_C����[f�J�������4y�~�e��-��q��TQ���Ql��a!\0=v�����$lp��p�	+P �r�UM�ߡ�����1���`\l��+q������XUlu_w�)�����K�(f�JG��+�EƆ@ga=���;�=*��2-��P��ř:j	�h6���]c�eDrp/N��Q�AH#�[�)�.Y�G�!2N��ۣ�~���9#�P5�`��[�Y>�E,��z$^��)�LM��rg[� r[V���Ee�n��W���tg���$�Z����m5)����o$���b��SPG����=�2�Z����≲T�2z������F��[$gU^��G(mERn2ѝ�'����J�7�C� L�G�N7��!�/��Vm��P�Ңp/���5P(���EJ��  B��%RW�c�38,��YE��������e��e�����\�ygO���:��oF= 3�O��~���@:Ez���/�z]�;>px�y�w���O��?��42�g-UT���tf�����s�O�{�n��FO1¡F�߄��wO�&Ԛ�gX2��MaMK��N��EEa#����(��eB,�s� �y��d~7Ͼc��a0�+[fG�fb�r��H��)�����,\��2�G��{�⏚��3�睰�͹H�܌}^g'ϝd��2���7������w�Z��ĵO ��Ω�h�~-=f��Ǯ��y��NU"��N�:L�_Q$�|�zN��jӍҺ�=���`���<�{�Dr0(��5���0% #���#�Dg�c�/_�m��`u�0i_�{2`���~��p͔}�s7	A��.�^è���#��f��W�~^:���o�4a��ϧu�ώc�B�p�P��'�-?�ac��x3�����,��E�ņ�����qM��޿���h5������H�܂�·�� 
x�z��,�t�<�`��N]��{�lϋ������p﹅b��E>M76ݹʷ��>�<o�R�X���~���K��'�z��� �ϊr��Uh���Ӝ�"�^��g�^�k�����b�ʫl���Ju;	h�O+}NY�l�3�Q��3����~�BL�S� p �p��S�>@�y�v�䑷d�^�Y0H88Y��8r�=�-@��Z-�N��7Gw�ћ���;y��� ��j���%�ʿ̓��ǌ�^��� �,���:�M�G\91�݁���׼���`]�gw"׎�@���N�'��1�١a�;�`.Zc�[�?j��Wj��?Y"�d��C �pK�܆a���1S�[ʴ�:��1�-��k�c��lN�u��}��a�4L�.��.T���{�9�{7�h�h�ƍu��\��=y��Q�5��ӣ�s��/�L��(���~1�T�h��6Lr� �Ш�J��^/�:���&Z���מ���Ƕ�ut���ۢ�˧t�/F���,2-�sF���pN���CV(s�gMȲ��_��1M�8{�]m��*X��,me�$���	�=�)����:Bk^�N��p�W֋��@���_s(gw0�2�R@�A�Ѯ!�$�;�jk)%\�UC�?p�$��e@��?ذ����j�8����?3�ϯN��i�G���ZL��s���
��QqN������o�\(��;���X �B�(�mA��"2�.���d���vJߦۛ�K'��^M.닦�YA��w�1!�7�7+~�}��������C��~���Bҁ[  � �����,taڰjτ8�O&}�b�.��ٕ��L&�R�j������A��?^2O8m*�Mt[D*!�yƀ9@,��\�������mۍ�@7�HDVM�`�6Μ�<�� ���r\}��U�� <��:C����c����W5�O�ߴk}k��4N�1-�c[7��<�����`/��q��� ����x�6>6	�~]�k\��N�{�e�Wx!bϟ�t^N��������������ImJ��!�CB�D�O��ul�ǭ�]�]����?#V�]X�@�#�oMx���+�(�8�1���	5oD'�9|���L�)����óm6(`�N�J[��+���⸅��V�����lkOhpZ6��j����
�'"9?�S�ub���'��ךZ�w}��ę�ވ����%����L��3����TZ��E���;'�쳭�lθ�%�X��Lᙋ[}�;��g01ñ�y5-����du�s����B���l����Pp��ƄG��$���>�]�M�\jaU�������kd����O�����c(����ǀ?��|��7�c��	Z@�;l"�k���v��&�h� )�rΆ��+'��/�jۛ�0��6�߷��8��$�J��#z�$��wB�f5TS%��"���/N��0+}�Jʇ���-P��8$�b���ԫ�����("C$�{��Jr�BO��   G �-W��÷rb�7��J�^��I�)t��ީQrG��[D�Ex���c7&�����>tEF�jM.0-۝9P_�܃��qM$9�n�o0��T[�"���k�2��~��Ϧ�hDD�"�`׌�L2M�HZA_|Id�� �sF���+D�SΆ���<1�;���Hwƺ���G*ߝu��&NbB���8~�)���~7+
�S`��'\+wX�c@��֜(�Шa���@�$ ���ݟ��?9���So�j�	�`k� G]��T8������)_[͊%7�1?���%k�Y��Nn߈��h<g~ 5�	Ǥ�q�dSky���	��V��f5V��؟��g�E��AΎp�3�!�����sǟ�hO �=	��(n1ş>�����㽁�=r3�Ir�K�H�;Ի��r������&W;�|d�����vbB�k��=�?��
a��o
b��̈,fCS\N�e�%����.����^W�e'P�|r�L7<�S�/�E��.�4�Z�pQC/0�e�l�k�!2!�����J��h�&�ǩZ�^V6�?�x:�o�P@��2�����EA�f��������!�▏ @ 
V]{-@ [���[�)NP�W�&�s�����"θ��Z��H�R}5P�q���t��*�'�S�R�y��RJ5z��_�Vm����EmAyZ�A
���K7j@��h7<������o˓���  �!��*��1 $1H��� '@,}���;2d0��C��?`nڻZ��%
��<�?G�� o8M�ݶ7�ݪ+wlճ�~�V��e�b�+��5>K���K+R*@�X*e�驆T����W����9��2�ɜ> ��C�k���C"�   �!��*�b@ �]�,��%�MȔs��g1����$��P�Rf�FS�u���G�F���.�$6T��!f�6�S����� �;�v}� W�ݧ��G�<;A����v[U�!�Bw�� � �5�@��@ ��N%8@x���[t�U,V�#��0  8!���D���D�ܨ��z
Z�,,,D�U�M ��W�Vy����4����u���h��9e]e�pw���I����
�ݷؾ���vm������/�B��d���n�����"(NR��~�����.����G�2�4��B�*�y��+�����m����cz��   �!���B�lN+�nT7`@D4,A`@��u�B@�����M˞��7.p0��iL�ۤ?���j-��7:����9����tE����+D� �r�aB]�C�TѰ��#�k��^H�"�K�2���. �B�܁Q�?�ߣ���WG�) n����xy�I���  �!���	B
B���2�Ya ��h-���@�N�j'��t�xG�(�1�g��7:��Aj[gq�*���s��1����Hu	��N�8"�,=�erD'U��K[05{D�K���zd�s�߉B馉�%�i������;����0/ ���D@@��&�{}:��T-Z���nR���  8!��̓�X�&B�R�j����y+v�]v��V�a(AE�O�J�Hp08�B�]��O�"P�FĈ�93���\�n,A/8ֱY����2F�#Yř�+�����k��i�=[e��9�D�Q*0��K��˟���z5x�I-�*r�k:L�( \@��F�ǃ��E��P� :6�l��}iۤ+�]���R��� �!��e���|�;P�P�@Y^/�R��8L�8��}�� �5��\�(��α1M��2����gB�u���ƾV�H�D�t�t�+�.1d�1�%�
_�Ǭ�?h+���⡼)�I�a����:��	�Xl�O�;���VS|���_�f�B `   ` 8�N���   ��p��W�C����hzp�KN�����c�zxQ��+�y������?u�1��&��r��!��W$�X2�	 yAʨؠ��wG�K6���(�Q(��U�8w�jm=Ԟ)�w>�T�������|k�98`�¾�$F���Ta1�����hKO�
jͤ������f@��tBJ\��5�	h���wa^nZ%[a<v��l�ٲ�lle�R�$�huc�����ge�bҫ�c3?'vz^����h�H��Ǩ�vW��ʡ���F]�dY�WR7���]s�ԇ_�y���:�d�AeE�ă6^,H�%L�qRd�Ӡ�1�ݟb��	���+��]~�n�?@t���cX��d�J#DK�/��6�H Rn�6d��"��[м4�����jc�q*��hss}��i�s�����y�,���D�1f�S��񀥌N��H��}9�<��2u�F�J�U�㤇&�?�k��b�K,�x]yD�J�����(2P~p*�H#d�����Q���`;��%���Z��%��.mY$�2���p�����j)T�f���r��<Ý��s�ȯ�*�6H�6�.C9��SY䡞.������=M0����G�y����xF���P~f^>�<�1�kO%����L��?�4h�a�}}&R��	0w�O#��"�渞�4B��p'�7�˵