m�u^૑�L�;�>
��J<DP��+-�)+�Ow�P�y��%��T�?ܚ�Kg�A��R�p��V�I�s�Ƅmg��=�h�9�04��m��7���R�9��b)�_�t��ob���#]`�a��&P�;��T��u��-�e��z����Z� Ô�.�6E����cB��+�ľ_
NtJM�9U,jlb	�����׀׀w��T3B\�]��Ac��T^���6&��x0Z�`����8�j�X�z|�+g���1򠍜ߤ�ʃra�c�.0��m����`��6k�B/��Hl�v��@��c�D5���<0j��\E�:2�
{]Ϳ��DIW&C/�1J��F�hs ��ͪs��ĕJr�E'����^%l*҆(l�@�M�/��ֶ�;��6~x�EY}f��x���ao���"��U�A�
n   � ���u�m�z[��7N2�_���ϴTAk~4�aDv�{[h�1TK�j��v�a."b��{�ވ��@���e�I"�FC�c-�'�.�jb���+���j3}�ZaұGQ�$�&&7->�u뉭$��Ǔ�������NK�r��l���Ù[��Add+Iu�\���{��Te�8|�����Ŕk<�Ѓ���赶���t�����I�0MkNB��r���f�U�����ԉ����"4��yy����>>�(��oݮ����U���j����
FJJ-9�I�ѓm~�T�7��;�CU����	w��-G ��6v���t��Tv
��j�Z�]7�x���E<@"�Wp%B��W��'�	JY�갬�I�7�ff��?�����ԩ��Á�TĈ3;��҆Z&���<��e&�{m�%���8�Y�5�"�J@�]��@������g�5ڋp#��I~ߖ"i�=�@ãA��
�   � �"-���æTt�J�ɖ
2�_�%���հs[�4����zK0�����8b-�V��MU�3��&�����MA�۾6�/��ԴF��\�$Z�����δAM�䘅��-k& 8����ǹ�������i�/��:g��P�p���hRp5��=gDzMǂW�(�c�
 �b��Y���ʔ.P�q9�����WB<+�G!�U
�)��ͫ���ʒ�K>��1�L�Q�W6�˗�UWr��\`�\LD1��R@�*�"�(������^].�Jn��m��	�!������C2P�p]�%�:���J�}y��8�%?.(t���y�r_&$��e��dғ0!U�m\:��#	� �/����}_ƄV��t9z]�:���{pm��y`�/��q�F�\/�<�E �f��������!��"�#�8�N+	Xd
���=��6�A'﹦�a�dJ� �3� ����5G+�M�h��`H���3�?Z��?��7�sw[?�i� �Q8���BA�_� '�a��s��� �����@�09`�?`���H�T$�N��A�HBc��>>_K�~� �� !��"Ą��,(+P� �T��)�A��6sS����&RW��� R�~j�ۓ���;������΂����@�7�l��j�<���D�S���cg�$% ��ˢ� �,�0B@0��0I�,f��� ���H\sv~^|�����  � !��"ă� �@*  5�~��A�+i�!��ٺ3�Lԉ�.=�G?_j��U)��툟h�q�N��i҅4���ێ�&E[���w����#n�h�(��R�)��z����15�x�`&Հ�H �нxl/q� 0D]�s0D�
Qz����q�w��   �!�
Ђ�l�1@	���Y�*PC�5��A�M�3���� D��d���[��;�nJDi�-��y>O�ۯ�$���G��e�q������7��6G󽿞'�3�C�h�p#V�`2ߡ^Vѣ��}�Bi
����P�[4���Hn�	}�  8!�
����@b�� ˛ɽ~s�/������S/\��0`�{}�5�@
'b��`:�M�(2>�^4Z�urv{���]��.%��v�l��̫0�J��bHB�(��\���v.MC� |{M���+9_�ߟ7���  �!���Bc�B�G1V*"�et����Ҏ�*�d�f!�X�+T���n�<f!��>� w���Y��eP���7�{~���L��y�u��I����K?�޸l!&LQ�����fn���z��>2�|�N�!ٰ�%�}x�`  !���ȡ�"�.��iL�A����7O�H��S�$�����uɘ��[F5���5��悥N]ڰ��$^?Ɵ�Ij��H��6X��� h*2+�k�,��%�7�W>��ze���׊@���<9[r���8!4��@�!��*���OԼ���  �!���ȁ��1y9�eI�kZ#jJnu\��(��r�c� `�h!ZAȤ�<�a"����Ò��S H���ܑ*�/�w�^v��U�����}��Ѱp:yU�~�Ϻ���H%�IU pp�2���\�8z>�4���%+��	�|���Q���5�~i�7��   8�KG��   ?�8����C���,�v��Kq�_�,���[ Mm�c�#�`g��b��ob~��J��Tv�`Zb��[;�l�@��Y���&���v�2��LNZ��w�]�:��m���޹�*�*�11C9ݟ��#<����#ȷQ�K�T(�,��y*��`P��C������-��;9S��ƒ��\	���!�V�����ج[e<��qɁ�'�X[�r�O5��(#���R���z��8>4�s!���� e�����9]�'�_��v����{�����~�q[�A0 g���~<�+U��Y$���6���1�ۛ�Tl)ep�x��۱�g N��|E�o^�[��ΐI���B�Z�.��rO���.#لX�'avz�S�����m�����RPD����=?�B�!�����ʑ룫��eyIx��/�-꺡�T�j.Nh$檎5RO_%��:�Xo�J�p��ph�d1�`�z���]_L�c��<A 6�8g
�.S�3���T��L�R�RA��]-�DPqy�\(�y�M'�F��<�W��&���Z��K��@h�A5d�n�hb�M���*P	vڿ5�����U)�X����'�8����������T���'�F���}���Xn�K��)�X�.��a�0H�o��G�ǃ$�U���npU�dXί���CxJƣI�>�
�[�V�|԰����jHvD|��:��$+C��/���pkg�l!�<i�l/;�ʉ��d�K��g��뮋��\��e��y<�J��L?���{�8�¼��]E?z�r�}�W��e���7�t@fV�b�ƈ���_�Z���KA��w�Ǡ�m�i$i�{���0lòT-�1�Qo���?+@�xp\h�Wr��-�-u(�]w�$- ����aU�beq~�dВ���]�T�)Dq��0����Wo$�;�q���;9P����t	^�G��W�3������OZ���|ixD����[�ʚ�K�'e��&AW'MB�-������'0�Ÿ[O�]�^c��oUT)me3<���