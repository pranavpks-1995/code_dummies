H�WxC�߹b�e���m+�h�sUg1� �Q2���0�P M�٪��Y�����ZF��)�:o]~���C��q'��
mCA@�1n�"�����*w3��t��]��i3�2�n�t�W����l�����S�#IRq:Fޡ�:��5�!e�<D�|�4/U���o�����u�d{OΕ!g�Z8��[p��*U�_�s\j��<!Yj���Cg�_�R�,����u�j�Ut�'��=�g���� �!�5B7�v���i�S^�:)4V�7�;�`ȳ��VByQ)z����`�YΡ@Ӌ�WR3>�������kC�#�!��5(�{����`�N���%��#ap�{�U�Ӻ���O**�H	'�3������[�?�\�'�`C-O���z��#�f.Y�E�*������򑆕�\2R�M1����L��@��f��ƪc
�����/��3MKu��\�m���!:��"�Q"hlF��䙅DU���Ca(O�y�Ȩ���0;���;ث��Z�r�m�᭸4;�D�`|���pY\��[��*��\ڊxĪ��-�<���̺���8!h���X45Vg1nOT���ߋs����P��i	�����+3}T�p�	u�%�f0�8`�"����_�:���Ab��Wj=k��Pt�!1`tά��±�9]0q��=��.�QI�{����~�F���}u2�j`d�� ��>��zc'H�\���ԗ�����l��8���c�M���)28e��N��a��n��$�� ���ӟ@$T��j����r_�f���T�Vu�cka�Kig]�Ñ�N��A�(�G��������^la�����+P��sR%5�`�51]�S2��@�����
)U����?M���S�.��z9�*2�h���Y?z��G��^�}�t'��,��)�(�De���]��_�|b�T�����
�(bdP2�����4���-|�
]Q��4w��#�!Tq��:
ΐ�4���Ľ���!�Hqh:���e���0�~槯�ɴ��P�����}�v��((�1��b�M4�.wu��^�g/��ֿ��rB��[�JVF�"���~A&���2��[u�1Yq4_�x�(�g��~�UUS0�.pO��9�H�"��z��z>�.���s��{�P��pfY
��Ld�8B8��z��J���ԎML��rY������$����)�u)n��	{��ͷ�a�q�.��E_E|�����,�q�N!(7�_I���g�d���Q/O��a_7]����¶����E�|@O3��vs�u��#���@4�w1�@�1�	I:�v���&X�}!�� ��?�+��Y��,�� V��@'�l���-8]����8V֦�/��+������D�HBbR�
��%Z�f�o�-a�U%#tԫ�
��h����8�Qf=وb�H�I�])����0,����d�"�9[��;=�#"�4J���������eetEpk����R�J�})M��zј�����d�{K�W ��g�Ρ�o��ӵ}E�Ƚ=$�n+��߱��A�g����@W��6R��i������j�{��4�0W)���虏!����r*�r���c�Q��1m��z9��]�k*B#�Qr-_���G� F�d/F��t0��P�N�p��Yޚ�XkAc��]��o��mȈD˝�EC�[�17N��R]�ԅ�8��|�`vTw��b�<v�&'q��#�Q0Phsr^��Ȗ�F"T5����Y��Wayٔ�B�t�GSdz*�8�w�a��4�d{�"-,
M� h�ƈ?Н�۪ ��f�M^�,�xW���F��IY�_qc(]ż�	E4/L�;a˽��9^^�r�ܽa�>���W�u��0X�G��v�pï�cӛ|i.�'��y:}m��E�`SB����$vޣq$���%����n�VL�I�!���/#CD	�`8M�"�F�N��џ�b�PL����Z@���Aq����T� ���?�`D�?�*�Kd��W�f��h��N4��}��l@�]�XV�� �L��zY�b�_��q�ѐ�r��Ƽ��ɒ�C����4H� V�&
u�J/`�����	]�.6BI�P���.Y�V6&�f��e=�3��\�>7�"xd�����i���J����Ę�_f`��B��}`/�uK����NxB�_�wro�P�䰊qeW���r{��(���)�T�
F"&��YgP��ڳzjȩ��㒸CMH6Zޮ?��J�����iB9�����|/�{/��|RczΟx����d#�v�^�E!�	Fr=n����H�����G�|���'�� ��U4�U�n��s�~(޷=αx6^�֟+渠���~?��>\�B�h`I�!~V�D�-��t�2���\r=�o�����������З�3�����c���q��ע�|�3;w�Շ�d���b2'���Ƿ����+�e���+_Pb2;7I;Q4P�\lh]�\��J�%�x�~��T�B����**��r=/�ݐ��/Q�՞4	�yT�o��Y�<NVO�!�E]M��$���T}��;釲z��J'Ӵ1.���o���4��}
��k�2{Q��HT���H+��)�m�����r&�g�F{4�<؆m�;�я�⛭�;-}|�]�=a�H���Ov��X��nQ��08�Pǉܠ��t�O��������|�ёb=�S��Ħ˥��e���Sѕ`�Z6���I�G�~C��F��k�<�x��m �3�%#O���[@�a cV!�ဤ��֌�a��k+��dfe�Έb�s��{��Ԃ�1PV�}�:�ܥ�k�� V5<,��M�m_5(���o��/^?`(;��Z�5�HFic*�QnC��rm���&=ԡ
=&��C�:���u����D�=�vv
������[D
BR�E���b?�7*��Ǩ+:e���1�M��z�^��@��2�pn��#x����A����P�t#��^2��<5����AI���Qc]�\���V�|�l��B%b��5�%�Z�n��i�4��p}ytWE�46��'�|;�~�����*繉?��+a����U��5�ph���pw��&�'v�$��ȿ���AY*o�ɩ�i�Ccgs�H,� ��8�Sb�z|Ӗ*[����)�n@M�L���j
1&�1'��R�̩x&������	���L��F,[F)�}��B�#��8��k���dC�� +r$؜�]�:��7�k�c����¾l�.f���BU��t�X������;a��\M��Z��ڊ>eԹcvm���Ѝv�m��4�'Td��Kď�݋�{R$9V��;�Q0O�cn�ѷl�#P%+5�����~-��@}G���GZK{\���"��ה\�ʍ�g��p
��\��)�}L���	���p�,	
1 #$��������#<��`-�YD��+�6l��Q8h���В'R��z�Ɋ�<��s@�;�-Ҭ�����W��-�a|��=��v��˲��O��*���Y�6ۜ��bF�/���'�x�9�å�2�A�\���Z�3?e㴡R�=슈1��a�v�� ~�1�r���:��z@W�-�;�X�F�J6��w&Eeo:�c��7������\�a�_~��ÿx� A��~j�����+u#Z�P��n��|p�0C�Bkn�8��$��{ֶ�Ae9�`5ϸx�G����n�\�g��:��ȳYv�e{���V� �E���  ���%RW�c���	U�`�6�$���Aa`�qaX9��.:䫭k�l�sKK:{/��0Λx��߿�}�t�����V�1��רu���xn�4ݓ#���ĔJWBش|=v�#̯ (�t �>��򡹶��<��_,����E�9�V��b������fVU��;zR�L��'�u;�� g���y��t��������H��@b��������"}�g�Y�n.Ĝ8G�'���Ε5��:�lҵ�����G�J��Qe5�������p<������(QF��:��ߔԇ�,l����Ȟ�F�$h����9v�T�Vŷ`��؇�(������g\�E_" ������vRh_З�29 3�ȏ�FY���x�Ԇ�)�.�V����~�*��LoZ�y/��}E�I��S�BX�y\h�"m�2�
#��ٸ������j�����)�C[���[D�����X��Ӈ������P�h�uxH��0���)I+-8�A��я���]�XtfC�������[���en�۴ �dF��-@������O7q[��=f�	&��vNdr�_�9�~�"�Õ��?��x3������n]"�-�H�w,�d���G�n�`�92�$m2�n�+C{�LN8@�E�RS�jk�܈1�6(G�L!�_�gR� Q��j�S����g��Zqy��8	�3F�v�;�gߺˠ�K`���"�p��à�X��"��`�Ð�<lEp}u���@��y�O��޴��sv��i����95���"�륞��v����W��H�|}�n�`���p����%6��D�
�#��@�=#S��q��t��[HזJh���C����ӣ+���v`�seDJ�e!g#1,����t��b>��2vS��C�����5�\ j�3}h�a�G�&0�kl�W�O<�{s�q4vwQw�ˠ����]���?]�d0��iu���1/�Q<OQ�k��|�p�Ӧ]�d���06{�ųaR ����\��kr�	9�z�=�'$��3=��n$��SZ��t96���~=����jw3f�C���Ft��GreE��9��f5��(�/^�9��P8W9�vt@�; a#LA��C�BW�p�p<��8c���jl.�6A�Ώ�OG�ΐ��8�;�j�ɘIW,��(���B~-u�&3Tx콑t��k��0�V�i���i:k����ay
'���e��)&���j�����M2�nE~��Of�oTg�5��(�R��=m�}������й�Ȍ�pJ}!\˼G�+An��a�:i�x��MD��o03��!�^��"$����LP3+�|t��<t���%����԰x[�%U���fg��"�
B\𯸱W��������!��,m�o�ץn��ˣBo�W  g ����,t`�cT�� �x��Aak1��ǵ�S����_oW?��7u �GN	��hI�h��Q���b12>L&32�>�Z�!-J��͖a�$=A�)p���# U��j5�=��%��ݽ��� �c���~dta�1M��4Æ��0#�Է˳5#�B~	0������	��£@�Q"س��3Ҍ7��Ʉ��W�0XEXk�ƝK�nW����S��<)�����M2n�{�����!.�TeY���c�h,A�Uc��=jй����#^��I�`�$¡,B��D���~��@%}{��8̻NSZv_X�hE�������M���
��b�|�nK\�Mw(���������5 ��Q"�j���V��_���n�[���i��5Q�kLc���lS�M;�O�!��m�����F�)+(��+��#���}��ǐq� �?M1�f�b�VƟ����h�������<y�����E[���]N����\�$�",��ki|�5��<�p�����F �)�����!�����	�&	[�D��Պ�� �� �ܝ-D���]�,��@�Z���,�m�� �W��xWX(ne�@��݃N�-���B���   � ��-W���
燌�F��C�����F��Zد{j���S
�Om�$j�^�ܴ�1���pR'��f���*N6��,�[��q���e�E�c���v����أ�^PV)̼v�J�s�䇾�"!9�T��
���5_~A�HCT�ĳѦ-�v��b�(#M5cQ��h7�Z��K3�غ8�3�*�=%���O��9D�������^�w�����������J�*4.�w�n�(����0���X�:
��xزr��� ����g�� ��&�|��Y��'o
9޲:������$p���"GOw�vG��!����d~�.���~8DX��������>��rsT���B�b��%.��0�K7�H���Ąu�=s�7p�Z���a������LX�����H�6�	��M �^�5���C���/ڿ�41iɛ�}M�[�`��7���	��:�=�%DC$�G^-4~�wЏ�5�@���Ǿ��<�3o� 囤 �(;�j��K����$��R��p9^O��28��H2 �|o8�D2g��ת��Cg9H>�<��_�h��~��C���.V:u��`+������n*�����Y��$@{5Ex�>��'�ʼ{�.�~9D.l�l������DB��΄
,n�!��[���   }�(��W�C��{ĴV˿T[����\�~��`n䟅����(m��d�}��&_��?��L����{���n���]�,OE��O��Z$B�w�U��G
�0��%&vyH�zW�)�Dzoz8��'¥KX�����NF�4$~H�0Z��UJ#0�B��̏-d�~��3��R��vt���*�n��6�f�k��6�´�<���/7�����W��5�E*�}�V���3���9����X�*��J;����zI�|4�Q��M����.���E��q���첇��7�r����6�1���Ek@ઙޫڢ5D�kbɛ�˕��O�&�f��uD�Ʉ��z�=h)͌�4[mM�
�q���D�6�-k�t�!G.x�A�>�,&p\f�T ��ي}���K���g=('q&X��ɩ�E��o���p�$!����r�ׄ����d&��6w˩���Y3��gP=21�#�����
)䊅���W��sY����V$]JO������,XI��F���P�2�������Mv8�$6sX�������N��3�/���|�qu$���X�y[�Ȓ��o�\T]��u�� +^��?�f*��0��j��թ2�s��K��0n�$*U�A8	(�,�Tx�0H��_ �U엇�����e��-�M���?�kI�zS'&�s�H*զP,^��>��ՙ�iv�ջ�\�t��I������A��zv�cإ�1���f����7���*�8�B�.hf؎�ʕxZSD���M��u:Y�_��z����������!�9n\X'45l�5�;0 �W�M�_ c���H5�(15p�,P�ECgI-J�POq�+g/a�L���nPgr6�"�Z�B�I��=X-�
xF�&g�y�t�?�E�n����.0&`$`�^T�#�*��%@͵Vx�j�����dl����+bVW�6�3�f��?��ה�A*#�t(�Jw�>N=_��S3*��% i�h�}��	S1=s�R9;���@G�W�5� j�4��-`N�d �y��vOѲŞ3倿=oOOs�\,&
̌�G�k�AJY(�������E�H�C�H���1�X1����d�7�)bk\)]ۻ۞9aZO���dw�q�`>��1������ͷm�B<=_������U�;�!#�W�-:�Y��_�;�+�*ճ��z�6x���{uA	cKx�
��Qv\>ӣrB5dđ�LcKL��?�H�x���()ó݇���K�F5��K;�b�#!���͛W	�w����kzaP
�����eL/+�XcvM�G�Fa�����3��q]� ���>����a�W�,9K�~�;��u:ď���|E�Ĉ:�O����s�h�Fm^�|p�G D���	׆�����]y��Z�X��r�S���`���nE�v�"A<0��{U'%-B۫=�(?q�?�)���_���34gL�a
��6��@��}����,�U-�(��^�� ���_���\%�����Ni��'�����Y��۶{�p%�\3,�P�>h[,a!�5�z2p�����p�9y��-��*��ޓ�R?q1P��5]�.l�~������6NEѐϋ�umkɲ��RZ~]��#�E�y��E
�"a6���E�7��a V�VE`�d�ip�����X�@}*�GKL�V��a�$���8����R�vH��-W*W �2lH ?  +s0:<9ʕi�s1����u����hs���� ��R߂�+�b_��9N�6 ʧUX����V��d�)B	���a/`��{
v���/C���� '�.{ݼUӵ�P�z��J�u���"���Ҕ�$��L�2)�����r�	!@9�QF���~���ؽ{$Gj
��l@�x0��pS�G<:r��-���	�`,�o�!�}`uƱ�b�Kn�U'���}�Q�#�,�S]I��P�X�
z�atN�蠲r1�@G�J���C�!;g��٫ j}X�`��E~�Sz�AE"�AW�BB���4��ڗU1����!*f�+h�Sw������
��z>������|ws���悁�~�����aP�ql&l�+T?<[�V�$�8�lO$f��e��q�+�)�f���?�Cϰ�^� ��O�������\!��SY��V!wի�����18�:ex@y)�GU��D����b��=�������2.� ?�3z��R)�[�8��^!¢%U���*7��By�㰝[/+j��:Dn���>w�����X�4&��d����3�a@�D����UwY���o7�Gb��P���Z�u��`��ͯA^3��4:k6��T�oN,cb1�?P��u���+qr�LN�Q���H�&`��c~w�p�����%7����νg�6`�``��m�iV񭎥�-����� в2�j�{mD�[h-��X<m克��JJ[����BE6�m�x�l�X���j{`���s��]3�';,��!���d]� �Wg���𺞷���'Vq9����ӝd�'��+dR�y�KJ{�4�z�w�&
�+�n&��<cFB�:堝P!���Y}��$�q�I�'�V9( ����lx-�}��L�\�@H���M�\���-L��[�B����*��2s�X��Y�"�
9���'rؾ��aN���xgi㜭����gj5B?����v�i�L�2s����Wb*�n����jDfT���|'W��$���0��� �2�rtF�@[npT��y
)n9d�TDOMW#��	�H�ҫ5��*�:E>�E���T��G�oJon̵t�����ga�(԰��"�4H	p�ߵ��V�RM'a����m�rp�b���A�)����xb���hRX�m�$"��A;.��Q��nK�L˓:%T}_8�A	n-�����t�ͦ,���}��VqZ"bRU ��e��z��M�qnC��� g	Mx�9\��S8rM�/����Sl�o�x�;~��n��J���{�\��"^#0���F���gFz��.��&v^
��	3"U$Y�����p˝���J���ݏp<��
=+��s:y�E�sF`��L��}ey!��H���j,���<�M������bL/d�@�^�!�4y5�kC����`�֎�R�\1�"�Q�N�o�����7�rO�H>�_�z����y��C��3n�
��Q��4�0I�=�������8�V<7����[�0Jr�!#�e�a A���Nv�D���Ө���#=��'Ra����Š��|��h�(����V7@	���B��[�E3#$�_v%s��x-a�c�w���U�ʵ�aȮ����������w��'U��AOI��I$K�DaDڮ&�<�8=-�w�V>���U�ʔ��s(��P쓥�7����ӽG��t�1$5G��1|���x���E&-��<��nU���:ʉ�.-H����1���QS:	�Me��n���=�����aa��M�8��1�HI	r��j����n(�vt�^e��	#�|#�fn�.���m���c�k3�E{7��_��g:' �TZ8��X�HI,n�J�Y��`Z�/�����7��i�mG��i���oQ���ǆ"y��x���6�����.��n�1N��-;�������agY?���Oβ`%�{�DK��Go�s�h�%�f3Ei��u��^|��x�vS%0�����\M�=�]�|��ǜ��H�4K���i��������+As>+�4q��ŧ��o��1F�_���Mh�Ԯl%+�bZ��[�φ�l�ƴ6�|�����u��#U����^�2�:��ʲ��霴q�cmS>cz��g�~(��3AqQ�:W(���u��I7��tp~��O#�4���6�}(�n��yf�z�j�\��j\:yaa������'_2�/���خ���x
|*��R���6ŷ����,�ԼA/Z�'�?a�G�ñ��!L�G�>���k�Ӧ��[�jT]H���.�M��do\���z������ �F����拲X��TE����4'ߠ ��Z�!�j�o�C� |S5l��c�j�	]E�豐�Bm��c���	��n��v��w��N[j,v ͒h�'��Kq5ȭ�W��fϽԌ2�s���`��_F���m��U���kD^�y�y\�u�N����Ū�7��3-]-	�U]"�{��?I����'�r0�w�l7�ی��f�{�2����t߼��F撈^��N����0��3���_��J��6�Эl��`�۶�BR���7�+�Xbr>t����:�����G�N̮���TP�� �~ԅ3T`��8���D���8G�	��n�(����}#3)�d� �sY����&M�9ԭ晷�����������!]���p}�?�46Rq�w�N�U�:���d)�0�آ���.t�Nt��_��,�O�sA�j�ᙋ4d}�{��1h���J���H	n�Y��X>�����/c�"ֿO�3���MIO]z(�ݼ�aXk��ׄ웇��stS56@�yj��=.�>�ª.���4�\�"vI�A��>�5v��5���a?�[�_�fy-m�}B���D�)
���L{GB��J���ʏ>�,����$P��4Q.�T���%�.��{]g�ǐR��i�\��0&9�F��%���y'��\n	��s�S8b�<�9���~�F��V�N�j 'vM���� �����Ȝ�f���Z�:�P��7���`W�{8��0L���n���I�d�w�/�?���]���=�]���F17���@`/m�aF�����ؖq~���0�.�1X���Ms�.�� �����/њ�����-�hb�Z�~M����i�A��Tt�\[��O_�AO"F�'*�?F=<�!5u���ix���$��"*�V�u��S.��Qx����ޏ6	��Xب�,�CV�G�fi�|�Y�	���r\�)�E�>_œ��d�ۅ@�-b���� U����O����5�� ���7���jj�+<<H�N�����K�D'�O{��E��-�Ȥ�J�tP�G1Ŧ����0�v�W��O��n �Nl{޸��𣑭�:Xź�{*@�Ο[�X�tT�� v���Z�ԀyW�?����{S��+�Zy6����
���BA]�
#���w}ϸG�.�8����-���=u�v�	.�ɴ_Bq~}�Z���6Wb�%t��N���j���[�\o?�(��_�M�q8�ih	&yz?'�@'*��Yn9xѢUv�]�������k���{	����s5����!���š�e_��Ё����z~�|�J)�e�J��,)G|�4l�%ֶ ��Q|��x&&� ��1��m�$`kb��o�o�y��E��n߀<�ݵ~�Y`�.:c	k�| �OS��m!��)�����D���E/��2�;KU���I���Bb8�؋�7��M$�U�h��	��b/����J��X�H:�W��k��б���/iw�{�����O Qp)H��p�\������?�Qw��<�ɫgV�P+��U&��v�<芰�,\�,郍�N�L�*�ʧ,����Ѽח��"��L�}�D0ѱ��k �zM]�TYf���9F6?Y����^7�X|�W���}��Ђ��*ȕ�\g�װ�
�@F��Np���2�Z��?ߞ�IzV���pi<��Cx�5���9������[�� ��!Ѡ�4��X<��j�C-gL��w�{�M=�{*��_��u@���6�&�
M"��L&}Lh�\�@��mcg���|��՘��Ո��h���Gڴ��2���<H's����_�#u�?�&�P���K$��p!'S���Q�ss��t=XO,-�%�d~�`����R����0ݲ;Df��,�A�a��i�W��7�QB���1�+���� �e�#������_'��'�Lu �Աf w3�7�5p=���ۄ���/M��4��I=��}��Z���
R�)�j<���?��h
c�u���N =��|0B�������p�o���f�
|' ��C���֮9�@���m����k)��Cڑ;�prS�dc.4yk�2/@�IFQ'�^�^�S�Z�ԏ�F�K�N���~|�Q.E�]X��5�8��.K��'�*����0�$��{��e��t��Ws0�V�E��F?Ȣ7�<"�h��"�U��HT�"M�������iw��3������c�`���=Dœ"q&�e��ѳ֮������;S���P��e#槜^O3�_H�
��%���,*�گ�d�-F-k� ޏ�-�Z>f*� '�z���{YÝUv�\��ꓕ��Z�&,�X�_`�'G�5��'�hҔ��e\�՘\��rI��~�L�%��S�JA}�+�h�>�J��m!��|�����꾲I	�B�Q%E��Y�#sZ��B(v ��Z6-�SiZΨ��x�c(� �w�A�u���m�GQ՘ҭ��qʊ��h@�D�<U�˴7p�j|*gR��#q�K�.���St���g�j�A�@�L��Ux����j���0��5�\�R(#�{tMo�^1wZӂ}����"�h;Dr6�y�)[���v��x�c\�Hd��HU�2֭�|�H+�;����&P���(�^a�"�h�p-�ɝ��2eb]l� �Q����w}��_x{	�YB��NgDN��⮹C���v/Q=�E��3Q�Ñ���#�.�Z��<���:|1�����8W�K�l��*����Ƀ�NEI���Љ]����V�w;+�?�������r�漬��;��F��>	�/Y�pny��%��d�ծ�OR�ίc������˝}�nE�x��}JӔ0�?����^1���}oaw�e?/-a�5G��??>�悼؋�NP���{�c?��/,�Yc�U?��fG��$Il$�D<�ی��V�!	�E��'��E{zގ3m�Y9r��x��i�����8t�G�Q  �b'RW�c��G�\�d�:��征���ԧl�
���}ڛ�x�i�9�C��+���;��$)=L���{�<�6O�ƚ���8����%d:e��;�
�I��/1�����#(-��H\��7D�q"6oѾv������Sh6,�֕)�)��eUBU�7�a'P�n/`�]��Gf���s+�-(@rc�5J�Aq�/�sQᲺ��2=&��05@���B`]!֟Q������SZ�����	u�'ܗb�{�'�>4i��Y%Z�Όf�b�����f�?�E.�@��x����?�O�	5�,�b��%�_�
�`�y������}�՞�]���4��r���G1ݖ7�9�M���a������>�#�{�����T�S�D8�G3��E���\c7�7ޏ��u�~
�X��o��9��F��ݒ*�)V��9y ��<z��> ��
�($�ȍd����Kpz[��d�}PO��cՃ[���bT��{A�(�.�R��wO�F���2Ki���nr�BuE#�X���6�\�R,�
��҈z��� �
��~��2�!i�?��D�˘��7X�-S:\�%�
)��ۓ��Ű���ܱD 
^_��b��I7���%-�p�.����p��!��LUd����Bz$6mSׇ��:��2�/0=��6��>,�~S[��x۽�oQ�C�|�tB�г���4`�gdO��V�^1<Ld8:�����|^�������Nb
���z��3B=8���m��%�4���\�W��v�5X��K�1���௝K"�	0��s!Y��Ӕ�΁(U4��ֱņҬ�J��o.l*v������I�����U��!f�7}�"3�2�$��H�DЉ|��=}
-J�+��t��C�6?����#(�\%(X}��ܲ��f���m�x�4����I;��.�/Ϥ�+~/�t��5����H��)	zt������p_�� A߷��?7GD_���4��N(�.��s��AN�R�LLb_�q
��*8 �M+����i�S7U�Jg��G@hzi.���2�`ͨ�KdysI�Xc܌����=_ʮٴ�#���