t���?KSe+}ɛq��*�q��䀌 �D��D���+�ه
uf�o�@���EDk~�C���C.���B�a��Cm`s~�f�RB5
e�aꨙ����R�G��(l��|;u��$����Z�Ogϋ���?�	����jϫ��`�y�aT�_�)]�2C@�23隧����"���-��k�8'n��|A��
0���`Q�h*���@A3�&��rs�p�\I�0�Ў��������G�c�W؄3n��`�aj_�ڒ*]��8�P�
�	
7�k�n�Q_�6�S�pWwC{�q&�e��"[xݙ����'���1���MQv.�u�S!�O)�7�iN�R9~��bn�r9**��ܤ�tK��ۈS�B��G+�	��;�n��kx��f9RCK� �=W�W�a��vx�]6"�j���t��g�!��w�l�4���0��+l<�0��d�%ǉM"�<�M��S�2�1�7}a~]x�������q�VF�4[0�׆6�L�{U0q�C���K{��Ǘ�./� "���H��e�ǲ%�>"g��/�"']x0lh�LZ!�c�T&3�z�ٝ�	�5ۦȌ�IV-�AcP6:�3��X�C�����:�̀ �I����co�`*��[�W�O)�=���FJU�N�)���^�j:�x�����27�{��c'l5���:�I�<A�-|&��g����7�n�=���ז/İ�"�O|S}��R_��2xy���E�\����1�I��6�2���#��]�ݳ�k�7�B.8�ň�l$�7�7t;a.�b�u�������oj�g<(A\����K��š7MrùD������u�f�I?�cjEq��==�w	��=��MI%C���ZIir9;ӯ��U\s�F�����p�=s\����ROb@��@���,)�΅�Ϻ�x�$�MrNf ����d�0�j�w��natnE2sD	��9�ص��i��]Z6ڿ�sF�;�PK[R��5xa�l�=b�%�3�[G�^�LQ�A�����5ڒ�U�9����H���]ĿI{k��S�{�lb��%OIV�f��K.����o;RHm�G�DH��?�X.g�����<
�f�����ea�|hB��Lf��cx��Oef���f��L�%��6=έ�&Õ9���#Pe���H�"����&-�o�+����S����_՝\(.�k��j�BL��k(_���b�Le�sV�kZ� ��Wa���f�kk���1��]����0��H�W��	Y���}d�S6_��!���7��ֳ��7�20�4^����l�"��=XY7���Lf�j��.��Ҙ�H�YGH�@M�L6
R}�Q�Q�F.B���Z�w[d.B3��)�C�&�U{�N����"; @���:5Je2���DS��`Ӊ���b�EV��ȋS}*R�-��@��apQE}0j�IQ�C�-E4�ƊsY�c����r�7W;O���yYf�[u�Y�(�>�[Hi>�T���𚙷�J�!g.�Icc��^��P��m��H�*dM�&w��Jk�( �c��%��$�J�Ւ�}$���`b�KbQ�N�e���d�� P��:F##��Õ���9�N���II���e�],��a�7���� ���'�J���ݿ׋8ͥ����%�����Ms�/t��q�N��C
vWA�}_l�I/n�����_��Q���f�j���S��d�:{���O��#,�ݗ�;I�Ku����_����aY���e��9�ro���@����J'���3�hv�Z������+@����ɞe�	��T��1���OM��H+���j�qwC��c�~��N2[��u�C��� �Q� ��\.��_�ߍ���ˮ��hnHpW �5���(���g<Tқ.(�a-���Z#����/�P��
�f�s!�=�N6-�׷�������	���<����7�:�4�����n����As�J�[?�����
��w!��B�{%n+�iA��u^��F�4�o�j(�T�os��f]~?ľ��۾x��Z�~����\� ���D�%�����p��m4��V7����! <���rY�mRP[MȞ*����E���`M���U��	��#�{�&��Y_VT�rv�