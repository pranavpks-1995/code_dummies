package tracking;
	module program (Empty);
	endmodule
endpackage