���g��������x�[2�':P�UY1xշ�H@�(h��D���	/����%4[��UJ�S\�S���h9��WF��%d=�����H;�7M�{A�� ��~%;`��`��K '�����!�m��q����l���ye��{b�Smq��K��M�ғ�^�3.�%��T��e8�!ņ��f~<5k�lRV�^l�����w\�TEqs^�&,�1�2�*��^2�;���^�rFV6��G�\��p-�Qס�/���19ez�{)0
=��xfB(N� 7�R�U�.��	�7�����v_:H���.ދ����O+�
@�"�U˯]c�E��N����$a��n��e�p�`�G��
�"��F�β�Ӑ�*��B�V䩎�)f����c���TΈ�)o	���LW��k��u��7 �X<!����l��{�깄o�]��q>�}W9�g�/e���(c.it�Ƨ�n�h�hO䀶��(�XL���)��:�����R�Wa��ҩ�,�6��t�Pb�b��t$��������Q�V*À(��ag.rp�~�-�7;0�b���նG��Fx�u(z��5��I�'�T��D���e�c�AÆ~�&�)C����uT�������W!C/�*8وH	;����k��p�.��^'�&O�v%Z#$P�QB3m����	PS�J��q��
�����S�[��^��z��TO"Z9�Ѧі�R��*�yL�X��v�})D�I���+T�GT �w�ވ\�+���s��E�B��8�(e�����4�)j�K�����ڬ��Od�]�4��pT�L�Kk�7F�3��ş���$�Af�MP�U��`�`���h��%w_F���+�˒���������v���e���9Q�"i3C��J��QP�'�