�p�&�m�1��R�6��2�%�0:��^��C�ld �&��ݣl��-��O�a��h�Cܕ�ڞh,ʕh�@(&����E��)������S�o�@)�H���Y7�$�'�P�5����'����<����@VD�|_��(.b�q����J��c�tH �1�-�z�6�� ۂ6?�-ߵ�eF>]Z1{gg0p +��㧠�j�����ou0��f�E��	Ŵ\���1�������u�¾e�\2K�%�"�8ݼ�=C��X��s3Z	�V,�6����>�oU�J?������X=�sJK�l����`��c��C�y�k����"w����]['��}Bq��_��E,�~օ�9�$0�{��k��p.���`��ӀU(�{7�۞8�M���Il��wt�Ur:�ds�k~�H�=�qu��C.��ə�$�Wd��8�-�N6c5�t�J�Nܯ7����B���  ���%�_q��98K��kC%3$�� �Қ��+oN����_X�UP�<fq���U�f3������;�×Z=�uW�*���"��6���ybC�U(ŖN��?Z��Kx��FW���2a4%�M�7��L�W�j���
��_#�a��}�>��9- ML��(��:��b�«�k�k���w�ъ�����uS��i~�i�@�����{��ͦRhh�v�� �`z	}͇�