QР�������y�V��ٰ����@)���-�5b,$#�:�>�u��f���p�����S"��e���t�D�vh��P8�\����@˵�y:X��*���0���I�����s��+^8<H���k$��e>�]> T�/�g�aĴ7GMPɅ����G��M�
�D�ҟ2��-�+�P���>�2]�!ea��襔e��yƈ捓WH(T�JZ㺥��.w M�4GFv���G�|�9�> G>묢#�p�,�@Ԛ�?�y%_���B�〖�5kx���pG�?I�ؕ29���(���]��x��m6Q��G@�������9�#k�zL�NI�ෙ���'��DӁf  ��'R��c�أ΂x�4(¡��	gL���7����X�aAM�%�4�4�q�A���I]AZ?�����Ay���W~��9����5to�g���	0����v:���.ek�ڊ1w vT����0�艬RNCތ��"�~���
�Zf�朩�O�g�-�^��R�'�
D_ij��;�M8�<C8궳����!�}%�GQhY���%Z�P}l{�=$��F�-�� 2Epz�ta�Vܛ�w�,�����tbW�-����l�˘A��{k'B)�5t�3	)��GG��3$\H�=R��"LK��^�_��Zi��R\��۟_f�< ����j0���d=X@�������Xeqs�φR'�\|y(;��~-�<R솮���F��F`(|��4���]�Ns:���>� �#�����!p?I�6�͸eIn9��ik5F�r�DE(tA��@
��tM<X��ͷ��"<]ۨ�k��͐���L`p��PØ��m��M������EX�a7����ܐ��m̼�?�/oz�z^�K�+��h.��ŜXɷ�υf+ٴ�PK���10T�ã�	E�)fu'��r���,ANC_qq�RW��s,�Ԏ����H?XF�+N�C���C�]����&gCWӥ�H�
g^~zN�߀�7(��������ج!��_6��V�g��u�A���1S%x��	�] ��Z�W5��LN��ʤ��q�_� �K�����{��jC��,&.��ӭ���D���s�}?c�� �L`�A<�1��QvSN�&�#l�K�e�;�ָ",v��=��#�K�:�ݷw.8<:���{m~=�ĵCJX��|~mi��1�̗0N��xؑd"I7�c%�TzҿdW<�@��tG�y�]�.�@|�V ��/�����	\��nw�w[I���[�̑a�P;_����[�<hȄ��|f�X"�o6ȈY��c�Y���Ӊ��¤]��ZҦ>�����<q����[U�[�B���yrEN����ۏ�Y�}�,
�g����Z�R�Lͣ�r��Pȑ�a���`�R�?G���py֒���ß,��P��x�V�Dp���2�'��4 ��<w�m�7�oE�y��$��$$l�ژ�a���4L���2��/�Ι�"�Wr��ҋ([��xU��Z��]D��f=�v��z13�K���j