N��]���O �c�L� ޛ��c ��E���QB�܋�&a�L-��a�m�oWl��	[�e��3��Wz�rDE9�L�.�vH1�h��㰷%FӝN���O+yxH��ȃ�S����Ll��W]�C�v"��"� !��Y��<����"!��m(��nC��?=�t�}7�G�!�M�F� ~锞���'j�ZA}�0��b�:�����d�m����ފ�¡R�*�~�~��3�hbX����J����ǐO�Q��ӹo�F(��{2cgT��y+D��bir	�z[S_|����3n�z�h��$�mLɂ`�!��~y�T�n��߫�cj�_���»1*v�iԘ���$������K�ķ��ʙ~��|v�(���kU�3�d�vi�
Vaɫ
�goW�[�G��5e�/ι�����!:��Z դ	n�:G=�]�@��l��(
S�+1�Z
�=�������V���x(�U3��g��$q9�#��W<A$*��_���m#��h�2����[F0?Q�w8��Y|�aA-'��H��=��]�GI�����B8�k����4�dFr�,!�t���z� r������WL��Է7���nj������u.�/bހ$C<�5<�A
Ζ�#���$2�q\�}|!����6т�����f�L�ˁ-��*z[��7�̓��,Em�e��g��X�)~�(ĀM�Bn�Jn�����N���5Oվ�f��0i�k�cB���t��VISX l��!�q>���Y��2�\C�/5��8�*BdtH|�n���Yҵ�"��?̢M<+�������;Z���nt����6�o��<[?�8�g�����X�̄m*nܿ���lD�;(/Vr�jғ��py3�����l~����I��lL|1��,��TQp5_�39�W�7���`u3��=�������(�
AЖRq�4�=�k����*��+cF�#�YD�2�C�[c�̪v��܁b,Þ|�� 5_j" @e�����J5I5 P��>S��>�~�k]l|�P�mL�@_���x����S�ɸ&����_Fᙛ(�C�K��{�4�[�4��J
����M�O���zA��7t�vE��A��T�L�����;�fL'+���PXw�X��1Ai����O����Ħ��{�f6ԋ����2��˭$��Rbʍ�>�rX��&�^��P1�iIg������/�6�c��"���8���[��/`h�j#��9��=��Y��P�<�uw�N+��#	�,��R�����s� ��&|8$��h%�h˪�
U40d�J��  
��%RW�c�>n�������R �#�T�(����F�C��ɴHx��;D��]
#�	2�үc�CmX��QrC�;@Wz:t��avS�f}M5��{����,,Y;����b������qDX���7id�>1Л�|Ix��;� ~;����D>a3�%\�)}&�empҪ-=S>��>|j����{�W��ϗ���m�9�DC_Bg�C$��TH�S�+��h�K.�N`]���a�X��(t���RF�E�.�Ju�Z(d�ѻ;���|ހ�h�)�Z,K����Cb��L;j�E��&�m��rP8Uu�T��n�y@�9)�!ķD����lFq����D���`s�kP���d�@'?��2g��n�B!=�㝪�nr'�c�;��EIi�^ߺk�3Йp&�L�/��~$�(��}9������}2���{�q�)�?�bX%���&`�u4�#}�S>�Z6�!غqvgI���~�Ոo^�ttp��,�������[-+GӍ(�y�鲑� ��8�L����@b�,�B�aYX��c�=����|�X	2T	Y �3�����<k�"�L���~�~u_�l�Ot�f�Y���v��^p�+rU��ɥX�Q:�/q_ch�I��ږOP�0��>2�/~�)���̏�:����;��"���>a�B���Ad�7�@��ͽr���{Rt�k`)��/��^,o���켴Й�gF��j�� %@�W�C5�g^���-Lѫ�֓����\e��^��XT�B*$p�T��Ҿ*$�� �#�j"O�`�d�8z����M�+˘��39cd0��v�yX����dz6�{4������m$ow�?�\E������V$���g�`0� �yl�a?) �x3�����$�$#Z/���okߣ�Hҧ�""��c�E:��^{bA���h<f���+R��������_��f��7;���+VŨ��N�"���	�����).nY�,;�#���v{�%Sd���'H=6��pgd�vy���F1�nWn���&;�ʘ�����0��K��>:ꁘ#�M�{t�h	:d���1Ɍ�`C���%���p�Ή���g��'�<T�� å�7��Ҥ�.�_A߬�q��q8Jx����%/�+���yĞ��Ȧ��+#�\ �� ��4�A�J�om_���i�,5O�{�G�)j�u1�|�
�P��<�x�BCWJB�9��i����,�� �����W҈�8�L�G-�� m&a��C�>I��|��F��I�R������Mx��Zd�;��ht}_B�WUi�3q�k#������G�o���@��S"`=Ȱ��T�����˕�q"�Ǽ�Q��3��%�j&e[�I��]�u��!�s�ߗ/�/����'(�� i��GuɳjwX �4����Hc�ˍ,�j�d_ar�>4�Ⱦ<0J�uΏ����71c�W9�����\�P�KxSӄ-�d���qL����ᧂ7�i��~��b��������|h��H������E�L5��^_����J��Ωc͢
�R����$8>�&�����u�?�C��d�!�gb��8�+<rO�Ґ�@x��c�������}o>jfJ](`Cv�ڱ�'����>�[��s�d|Z�-a��_+���Ьa��#���X�~���Lb��d�R��I�3zV�������h��p�y'{�a�Y%16C�tHI2�`�[a�E�����<3>��^�V��&���#�$��a��iס�Pg��!n�v��`R��*���(U�ߟ�#� ��'*��}'��V@�Fԛ�N��W������,�
ݶGcK����Ƙ��)��(`� ]���r��a� 6m���w��A��_���M�,0�C�w%&o�S�����}���1<�B�� ᶓ^�jZN��2nEܥ���ͭၖ�ˬs#�\ӂ���>�����K^}�P�H3�����;NǞ��mu�1���wV�-�2�ha�X��W��e	��ن�][@o�����*ID��e�A�͖q���ޥR��i�}>$���oڵ�n��iO'�OZ����4��P ��ؕ�S}�A
v�}K^\[���<��JY��o��hϤ�C#�4�f�7Zg�v�W��\�ar5�}���_�]�jh�ڼH'ƿ�.�(��w����Z���-2�e�ǝp*�sd��K�$��ԕb��Hb%�<��r
Ǖa}?m
CoEA]kΗ��僻F"0�����n��m+�Eb���,M��,��h~�w8��쫔�EC߿|R�+Q�&Ű���2�=!��cׁ�� ���c`Ӱ�Z�Or�Upg�(S�5��7)�U@H��T�֠>������}ү��s��g��@�s��<1"�}����4[/�Wd\�����
;��d��M��_5>A�S!��}�&���`}"V*k˳�� _������CrU+�g�	"�G{�hX�Ev�[�ÊJ��X��p�%�׬����;u��?���k�� c/]F����\���V���d�d��50�k�7gX_���R��DD	P�"��z����*G\C
�P���h>/QO�3=p_��k�|�eqWr��:W`hY�Uq�%dҙ#࿓�� u{&����!�XQv�A�t�ef�B+�-�H	�����o��(����F}��>��\��v-�Yת����G��!�ͪ� GGq$􋡏�A��bw뺆�y��b*�E�* ��9ڙ4L���c�Z~��H���E?�a  7 �f���,t`��̾A(@�,�D��NI�;f|�w	���)P��~f��>k�n�^���� L�g���ℑ���?��iiχ�i�F���MH^��6fN�yBM6g�+��`�����)�-�4h�w�#}���/�>�
�$Q/U�U�&~,�ũ�}#'v� �V%�>���Ó���A�l�=p�rb�Ԇ*��v��ro�4�(ۇ�v+k X�v�Z����KZ%�L�������M5@?��Y����0@K�-P	&����I������<9td�aT{.��d_�A��<�"�X+��qe� ��W<v��"��u�T�إ�N}A�\_� h�*[@|�XP־	�J˶�z��� v�t���NlaC@�՟m~^���6����*vDl|N����	���0Z�C},%ay���Jô�l2P�+��y���$=�K]���DL)-o�[e�������)a�\��L��z��jU�y�Ӥ�0�3Z�����n��IP��0��t�_`̳t =e��t��G\i[�o�K-��� ^W�+>AܝN:���!v_kl�$R�І��
>(�G�3ȯJ4H#�e��줧�B�3����� �uï�c�A�3�c.袵c�  ����-��yq���C\��)��9t� ��s'��䊬�8��^�y�����/�bx̮�q��a�82����b)tql�0Gd%<����m{5j~�S��|�#�dܱ�U��7"Js�Q��ś�B/w�g���[�j�N�PlRɹ*ؐmy�+�_BV��c
�`��A�q��~�I�w&����4K,j������@��y�(�!��N��;�&��o���Hm��ⓒ�鈝���Jh���D�����Zkr�~�=��㠹�|*JL=o��	��EX��^�>�"��efJ�,NC��_�~�e6eh�=w�Q�ԕ���L�ĉ�ZK�`���{dH�7d�?~μ|^��xu>�x�s����������~H1lq�*m�G��t��0n8�!.A��o��ʥ��Z~��Y����LIW\�zY�%`!,JRN�.&�;FN���42����߽��߯���jL��t��g����+8�������Z{�4,2��V'E������G0���z��!���rٶH3`�~5�D1�?���A�R�am�Z$�[2����=D.�!�2g�J{i������r^�$՛8�+�gպ*I�U�ǐ�w��^�/"�Fm|p��*6.��am�M[=Z�_�)�Ș�.����\�y����5�iA#lw%���Sm���d@���{p�DY'��Y`  ����]�ay8 �EL��   D �-W���-���rkE��`V�E�+}�X��6=����ޭ���|��Ȥ�R��"�n
p�l��/�e'{�luP��J�� ���i�@�O+����Z���B�W�]`���L:���.;7)wH]���s���f��~��6m��L!��*�F��zL�ۢj(��8��!D�/�`U��[��Cv��1VH��5k2��Ϧt�Zsۦ�ǉ$��u��{�l��/�XuA8"B��@T��d�v�����h��2�M�YN��gU/�5�]%�So�o9��km�ٗ<U@�Y"�JA	]Y��E��$��>�g�m|a��$���N|�4]���`������L9��
��ΐ.ō�������D������%Z+���l�	] X �
h^r\��\��R	 �F��#6j����޴�;��y2i���1g98؁�@�\(�*D���Y��2۫2�
��;���ġB=B����YUq��u�"���� ��.G9�Π��75n8�Unr3%+�"��z�Z�#x6��~�q�H���8ƀ�,%9.">�������@H)Ǡz���Ĳ'Nۖ?S�b䭱��9�f��-�Uf�}�@�&�]��"vt�%c�|�2�xkfS@�R������q��^�.
��� Ѐ���IY����֯��ݿ������л?�w�6�T�qO�����0���j�Pv.x�h������9���y7ɦ��&�M�[&W�$� ���^e/�V �P�v|��]5Rp�Ɯq��F�{̊���7)8�A$�,9� ���6y.J���Ƭ����J��6�2����ɯ�x���ra|���?S��kߤb�L15N�/�W*�x��@���`�#�:�p���<����h�$��<�����������}:����ŷ��v�f����|�s�Y���~����H׹K2'@�I��a-�@�KP�g�k{_ Z���,ԐS,fO�M&�s�,1��C��4�R@�,�ja���j��ğ���#�\P;��z�x�׫qp�#X�����K�1t���@N�7i�n��\Q�a�U�V6E,^��x�4|�+�a7�uN�PFe���&�Q��&@�=�\�����u	 `��D�ψ<�����vJX�8x���qĈ*`�R�dlfX�\k׮����QC���=}�S��I�įP�c���"�$�gq�2jS�	��x��B�wwz���P+\�oM���u�Pj1/��Ŏ�i2V��ۏ�(����!��Ǧ��W�9�[\��|�~#
�ͤ0��G��x�Ҡ�d3�K�2�Lކ�P)��#�'�v�? ܏l�k��Հ�c���   #�ѐ�UW�C��bf�S���ԥNnq���hт�~U�У��H�a�������*�>��&(���-��(}��:A\�>m�
��3����Z�,�ǉ�x�a����ި�� ����\ p��������ô�*�\3�|[D"C��H���g��C����:���r;�i[ǈ21Z��M����2=�V:��L��V*z�S�C<�o3&�\M{���;�\�� ���@3��~Y��>��5��d$r�#�Y�e������<�{������|b�v{P����J+L��"KQ�a�-��3��<S�^�%�����Vt�CVB�30%�.�CLC� Р��;R�P�x�+Js�>Bm�w3����F���p��(CR�A8HS�ü���O��QFj�Xٌ��;�.�~0� �n�j'�m|�nvWR_���G(�v�e'^������Y(t��2�2OQ������Zj#��2FM�0���}H'��`���D#B�=�F�l�m�1���(�M�Tq�1��v��H�*�$r>�7n�P�G+�v� ?k-���*J�����<C)�־x:=��GL�C}QR'?cư�Ʀ��梐�pKi�w���d��;Ă��h֮0�l�S��҅_�l���&W�cj�ݕ��4���G̏�BNy�y��b�I�)$'���=�*tfRok3�ȫ؈�:5T�<�-�f�o�d֔o�_uCQ?Y���������}���u��+�a��_^�+f��$\ �W���`һ^.81?}�9a����:,(��w�=}�m�h$Az�25����a��ţYr)��=N�~��oF9Ջ�1��쪸������9fA�.����H#�-��ӱ|E��#x��[}��1�:\�R�[B�+*�(�>��J���H�en����?��P��;�%�U�dy�uT��ؑoE�0�k�e���/��Im�@��z��_���yr}v�HKj�a<��[��=^�� �t\ç�K�؞y�-��<��I�@�]敘 ji�,����P�6����#�EF�^�� ;6�&
N���~����g(f�# ���㖕#-�p�%�I��X=��*��,�Q�� �<y�:�&��]RC]y�X�j3Eu���L����=�d#���^=��(�l��,R��sZ^����%,����XY�Q�7�%�s�w-�P�$7��u�1�!G�Q�dHC^V+��r�|�$(!6��'��o'��r�6���y��[+�F�	U�k�E�4�S��Qu�(���Z��r��
���p�]n2YU��Gt]�z
����|���S�	�O0]P|�x������mm-���|B�ݫ���8"I�"�n��Z�C��]ͭ*T�R�W;�	��ڒ�X�Ҫ�^�p}ve�E`�\�HTȍ��\��Z�^X��T�@�<�&]{�CѬ��xm�8�s"�G�w�<#8�@�^�ٿ�j�I�CM��7M��[ݨ�+i�E,���#7P��5�y��l��hTR�C½���{�U��g�� 0lrE�ER�n��}6k�i���m�T���f�O�o�w�6߉���p�nƿ��Xa�\�|Mj�z� O��c�_�H@�i��|�/UF��ɞ���&�(���&�����,�9=�Xq:Lm=�塧x=(v����ez�@s��`<l �l��Gl��$)h�ln
�t$�<�:���4�����<���ݓ��[�yR ��d��^�)A6}x��� �ڳ�
�v����{�h�<�w���`�S��>������"MH��Y1@5eT�\{��r*_6��B�|Ж8�@]�KhT���gl�q�{�D�D�/M�7��ݥ�Ş�cd�ࣹ�W�^)1��궖�ի�֓�k�t$���/��.D?���v\M�$���ܻK�[Y�"��"�o0�P�9��b�t=9��v��rIO��џ�U!�r?J!ꔤ{��F�ٹr��NHld�h76>��g&�q>����w��E��� ��ڽ���M��VIr݄x�"�2X�@�m�V��m"i�x;"$�%jk6�WSsS��1&�b@�+�}�;9�2�wW#c����y!��d u=��ŉ�l�X�� L����L^����@�n����:�d�D�*�/
F8@���k \�|��LP�