�mq����3�3�wF>�};��|=� z�:�e ec�ryrĠ��QZ�w�8�k(*�1�r϶��NI :����'�0%�|�Fqٲ�0=�
���`C�bi4@O~y����7=&qs��}{��R�Wm�n�v�� Ӳ�vC��p���{��&.�.�������j��a��Ph?�@�(��v��f�ȹ'@$'vR�k��cH�����۞\x�����"|'�y ���7}L�J}��? ڛ�>�X[��Zt'S��s�EblN���hFc�L��:c]\�si(|�?{1�%�x;��u�*�\��
����U�"� 	�Ǒ��:�E�V�?E�Eɮ�]b����"M豈ش�nU<�~�pB�s�޻e��N_M�O?�`�52��\N4m�jn`��	�ɝ�;����+�F�I4߸��95,�ǭ�	�9HnX"j� �}�%��F�{rqD٤�/���%�ʠ-�+O宸����A7!���ruǨA���*��
�2|"�\l,':+�h�3�5'��@��#6l8b������D�� @� _��o ��@Y�*�|`�����繴j�"����rC�{�BP�G�@\>�JVZ�!�T�M��9 �R@��rmϖQ0]��#�!y�3�>�K��l�,/�)�Y�-'���^;oW��d��k�,q�6�W��_���2�����C�!��:v�����n��'��QN�,q�9L�he��b�(0��EV�A �d��,���Kl��h+���<$����C)E �h��-���W���9x�s�-sm^�N'�5M���:�}V6�lu��7p��B���
����o�*��Y��h�|�G��*P��>����D��f%�Gb	��3�%��{Z:o�vb�J2�
!'q���g�����Uh�h��r�t�0�Ny��糝�L���ٓAW�Z�~���,bcgM�f}�S��� ����U�'�f�9�U:���R)������i�Yj���� c�ϩQښrs`օ3�'ƿ���?�.	u��lv�ޚ�d.�S6vX}t:�;m���D�R�7=��-�v�1y#�(���4WR�7ߌ�^��j6��1+�������?�T�+�q�6=8w�����̠]�����I�>�[T�
���Y[��hjI�%���*؄�?_ȁ'���o�x���e�"4�݅��c�1����+#�#9c��Bf�M��<���	�w�ߠ��m$j�,���w(�z������l���:AKk�o$�x��g��R�9���QQ5��9�w�xk6��i?�ذ��K"Zm�'��ԏ~��~���6#cc�.�@\Ҹ#�%�e�MFO��"*��\>`#q��U�;�^��H�삠m���NS��ɟD��RA���im�8�RQtE��ݕ7⟢�[�{��:C���bq4��˻lU��@�!d�.D������e���Jx0ٲK���P�����έ�a��]��,�T�s��,�ք���d�[� ��A;Ȫq�O�0u�F��@�\�$�/5��io�E�����.���g���C(~!ߎJ1�P��w�eEaWߓf;k���[[E�'��@�T����邜g��h+9���!�t�BcY@�i>|F��c�eH�nS�Dw��<-�^��򎛼�r���|�q:����x���&�h��ȕ�7���&H��$��k�޻ 	t�é���dm3r~��{z���2Q���̞����]yq�W���$2�)����z��K�'L�
={�h�@�z�-�Z7�}��I�`��^�ՕX�+�|/cdg^�`�Qr�f��F���?�?zyVjb�Z�[<r+]%�Z ��+4/�B�/��
c�j�t)n�у���m܏���3���:�d�����x���H�E椶��o�n��:�R�B:�ؽ'/_Q�����FV��� ��L˗0s�ɼАoYY�Xb�l@����9Mn$���j���C����ۇ"�8�o�`>�:S�C%o�I�|a�ĶN��y�4ހE�9�=�|�>0�k�"�1��z3�[�K��&Md�,�U����Pe-�2YXŲ-(l��+�ׇ刺�����������QZ����B��	J  ��"%R��c�ͤ�/��P��!S �F-Oz���?��"ժo�&6�@��N�w���Ma"'�R������@�7��Lx��9�V�����)pVk�jVR6^<[םCK}�x��P�M��!/��(�^,04(BS�U)4�N/v/�ݍe-�X`"�\�	:x��ƶ���������O,"�^N�?|�_�F�/d�S��8��y�:��B�) �L��K��`�&/�,���tU��W�g��r*���[�~�V��]��l�E0Y�v�ۼw���V�Xp�~$��� ���?�J�t�����Ih,A�6��b���=���a�q�������C��Q:�Ƅ	��)�u1N" ����ʪD5k����p��<)'��R��EQK��DbU@�F��#��������� &��y�S��l=^����M�C�(Dp1���u���
<��ـ�d�1��Z��a��*����
�]r3E�|�,���.��n��������X�@��Uy~]��"1-'w<�W�)�o�����m|H�̳)�t	�!�8��J]���xD\�ȕ�͚M�AP7�/�.b�S�{��7�38z�q.@Z�*G�8[T�"����AM`l�|�`�clf(���R�n�C��{�8��A�	    ����,ta�NڑsO4x�hQ�W�;�~���{�����󫐂o����g��w�L�X�]~�Z�&�l�6%;�@o�Ѱ�@������V���(GS>�$�/��Puw=c��,�P� (FЍ��[���Q���h���!�{�I�kԮ󄤬+Y�~���P��R�Vz��e��=|�]d�XH=�(��_r�
�IP�`�k^�gi��P�+e`XE1`�	^�KHeNfo��a�%�C)��r�-T¦�H1�&�D@8��n4y2A�6�1~��@��	s    � �B-W���Ǹ��1*�u0\a��I����	Ei�[�7]-�jl86��,\��/�h�P\�ȃ���}4t��(	��Y)WN�O���	{:e��1��KC�R��hP����.�G�����f�v�[� ��c���g�Ũ#^��c�d�m�$*sP~�"�%W�B�%����f� ������p�����1�'5`AjUM���E�������@��5'O*��6R=b�n�tg�?��G��
n   �Ԁ��W�C���a?ً�L�'`�Hz�,֓���{� 0RĥY�Y�h���Ej��=��s!\�q�Q���蹷�;�����˿{���e֗R�o�R���4�����H1�Z�oZ>U&�DHw���F��#��T��&�æ�#�{$w��q����[�^JM�b����#+��sM�=��ԇ���Z�jr�'� �[�у�����[�I��|Ji���-$�S��[F����($��K}��}��H�$,�����]�R��1�M=U��R���sPs�!m#�	�S)�ԅ��8��N_�2�0�Y�, �(�����a�jvsv��B��/�|�.r�Ul��H�Z��^��Z�L�m`Ru��w2/Kj�QO.X)M���F9f��$Q��
�*v��%*3�
�@&�Ǧ`QV��P`E�!���Z&'�S�VFq��U ��47���nس��¤���N��0g�����y��(��#���5Q���c΄@�1s��#�W�/��N���|'&yJe(y�ɨ7�9������0KbY�ȟ���Z�(^��o���bR$��T�[kC�
�)H��/{�
~��g���sL�(�=�j.��J��