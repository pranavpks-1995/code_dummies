W�r��}�q��Ĉ���Hx��z6�����c_z
��G5O}\�UUS�M��Τ+�d��?�	��B�`�j�?��^ZB� ��_ף�-L VQTuRf� E>q���6q+��7^��h���kT��L��5w��Y9eڝ�b�7�"��~��*_Je���1ϒ�I��Fp�,��D���@��^q��p��n�
[�#�O�s�cE��'�Ѝ[%2*�n^�O���6,�sR�<�F�����Y��#2�ԧ�cq�	=螑���|���J�C���(V���Dlvb���S/�U������Dd:�[�F�
�F�� �u���0��$,�~��b��\���㸣+>1��a�F�=aߢ��|��bn�ొ@䭦I�UM��5��B�zt����j/{�E��9�IB�kk�̤������S��5�:�̎r��)yO�P#��$����j�'?��G;A�'���NU_��o"��٩6
əϤ��1��b�g�����_2{�=2�$(�"�垊��
���˿U��x��=��#����J����P}���jһN��I\��?����P�G���Y_{p'�u��-h@�M0�rCKs�������W�7w7"�:��'�]r^��"t�5��p���7/�������5��ۼ^��8ݒ���J �Z���!�� �2%���P�{��=��I��x�x��i=M��ѭ��e��a�ߡ��	i=�g%��gb��!��h���g� ���S<
E�>�n1��t�a�D����@�p���� s����D>ĎS�jF¤�I?�s�W���?�@����^{��_Ldn��4FM~ӊ�`�j�IQ�N3��e���/ F��R+���^����r��Y3l8/��ۦ)q��5^nԊ�T�`����ؐv�r�L��?_��� �͋�q���`�i��l��e��%�W�0���wE@)�]T>��T���"�����pw��\��c+��4���r���^,T��'\��,#�dJ�~�v4��I�Hff�H���b�VIL�p\�p7��{�/~��3#k�F�L�%,Ƅii�t�ʖ�R��+�s�g���U!lF�P��,|痽� r�P[���_<�4�Ԑc����EI�v�g�$�,�M�0�T�(�d�ҥ{r5|��4���_~b�x��|�Ā�C]�<  U�"%Rq���μr���d(�,ܖ!+V��\%>�d�G��]
�r��Kk�\R�B��ȯ˒4��_�����l���i��� �<d�m��r��}�{�d�2�Ċ�.��}�z�#O�4�
�y�O��BzT�2
�;\ X�+=J�֝��q��Pe�t����_%4y}7���������g���xe��!n� �� #�6xFc��	��/Nܱdw�����1�L����H��*�.�T��}[�	��7e��ZR�10S=Ui����cB�R��`4"a��WY|��
��Y�v�N-���ݎu�v��G3�<U�[{Ƚ@b*��� �S�ڒƜ7��'��X9��/�Mz�	((���ߋ���rr ��,�WR_z��
_?>��*�9��Z->�5�$��nrl���J��3K���T�m��%���[3g.�i��t,�)�6�ܿ��y���> $<�)l��)2ݕU�s��o$����� "�Uن&a(S6�E�W�oKֺt��I\�K�ӊ��%lx���}�����4�I0XT��ٝ�C���n`	�g-�8���B!����f&
P�Nj�����LI=���(7�52�U����Ŧm}-<r�/� �_ ����! ��U���C3FA���^�=��ũ�VT�݁*(�H�^;l�b24#2~�&�H�>�k��Z�tM��n-�8O�(|*(U���ǋ�(N���8�1Wg�m��h@I���m��DEl��N�[YX��?�����������^;�@�l-�	�_��*��T-�ȩ,�fa���}�`�Yc�wb7��K!W&�������b�C�   ���H�ч�f\�Q�pP0D���j��tq�t!sL��oe��á~���H�x�݀��S�Gׇ'�`�,���j�.�S/�4�
8tuiX#"Lܵ�X�x�㫁��0(n�	v~l~��3Z\�������|OE���#ɲb_,��+,���fez��E5��^dp����T��p�|2�Ǔ�m�Q(���X`�fG]� ��9n��^Z#��ȿy`��gf.�K�;��u p�
�:�xI��p�'����h���M���vg1c�Ij�7�W�Y"JC�����­&��~�*"�7m ��i�5���VLf�@�3��������M�Ce�>#��Q�N ᳀Op��/4/��Hy���+Ta*�p���? uwm�>qߠIR��4�������ʢ�{��D_6D�a��D%(Y������`�Gs�.�G.�@��O��w,�R��ZΗ�/Q�	�\Q��5&C6�Ъ���F�+�4���\�A�h���uN|�M�&�O$��#*,*���	��ą�W7��]�_�V)
��E0y��Аhu�s|M�8r`�Z����*��v颮)z%i{W0J,Qո����ܟ�x����ǻ��7��\���/��Qx���K�Cfei���Z�.��I�}�J���������#�H�IO\WT���ȝ�1��;ޝ����K=a��C��yf�5�k���	F�9~�/������_��ތ���=؃6$)���Z�VcWBl7-��w۵.��
Ӕ?i������8�[�6   �8��_q:0\��-�w�d>�!¶�I���h���՟�ؖf�"�;�"���/�=��������2}HFXޏ�������4M��!E[������b+2pF%W-�q�8~�ެa�H��Ҭ%�l�ؐk5������ʬB#*�$��Dt�L��o��S���u8�`��nة=�YE+YB��wOP��i�'�p��:_����#͝|u��/(��qY�X�wNMʺV�g�s㝆y���Q$���`�kC��7
meL�)��n!0�IΆJD�OdE��+���;��4��m;�`Zi��6ꈆ}��^�����JF�}�����Ƣ�z9��+��bO��&:%8-�>\67�I�����%������T�����4KsD��ao���倾;���y�nV0b���R���vI�U2kl���8�M�o�}����-���QTÖ�A�f���Й�"S�ٸ­����t�Y�v?������?0NF� �uzΤ�|c+R�W)��Uit�eM*����#��� *��$�̆dO�+�Z'�����'��n`���=����|U�H�^#'�00P��%(Z��o��j��SisQ�r"f� �&1�8����`�X�BK�����2Z����9���X��2GO&E;O���1N��kO��Sue�:5`��r��8|�^!g :�&I��H��C&`1B���.z�|{2��'��~hk(ggG�>D�c+m����ʞdG��-k'����(T]�ݐ��T���Ʀi���(۴�{B��4C'Ç^��el?����9����Fs���!!����v�l���!i�l.*��xˉ�@%L�Pn�O�q�bVr�'��.�p�O�%4��U��D�Q\�*��K��<r��d���q-|���|�?+R�J���97/msz�HƜ��#11pg>6vؕҾc�	4�Om4sA�P�x_�:[ po��+
(:�貯�tX�&�s'��/��:�>8��-$��!���j9guU��ү �L��:��,2�x�I�jѡ�T��A���_h�͓��ܕ�'co� � ��(��<D`lIE���� ƛ�g��I�@Hd�ήP��U�6T.=�Y�[�`C�,��
$�(���#i�)�X?5�������!�t���Z�M˻(��� \Un8b���̽�<�RN����L����q࢈E�ɔ.x;� >8K,�s��'�|�l�Z�V�b�S�v��|����	��]�=g,�E�I��i�����9]9h�^Sg��i/��oE���:Z���9�w��m�dΏ���(��t�ۛ�= m��!oeƢ��uO\�#Ԡbe[�è�R2=H�j�\��Y�����n��NF訇ay�*��*";���h��������JN����Z�����A�#�J.�P�uf�jr��Lp����-�1ۼ�$�a��9o`�UOy���'����%&���z�~mg�:|���ͻLں�i ��>�D-Ma!����.��G5H�)C
9�M�jr�.�@Yu㎅���tϚrǾ���\�([���t�J�糇����\�`�P���B��w��8i-
�W�f-Q��<�,$%3� �#�oK�A"=+�j�������	ݓ���X*up�m+;dFɨc6%�[�Y��d��2U�,�iК4]݌����ӌ���0M�M�}��Jt�:S�%�L�4)_>_�Jqx�#�6����,>�%j����-��,H ��a���s�4,(�/̷Zʴ ����G
�d��+矘9�jֈV"����Fc^��"�y��.�j�X]]���>N�=7� Ϻ(ځ7#υ�`�2]ht<z�D�Q�ڛ�&�*(�c��7��3�d`EΌ:A�jp�ɛ���oDzk������ �3�b�y������r��-���2B���� |Y����w���u!��{�>�ɱ��$��&:�y]��,���
.p�,���b��S�g�Ā�"�;_�-�y��c�ϪO^!6��$_��A$<Y�6B?N��`l8+�5XX�=?�j���MUܾe�U