package Adder_IFC;

interface Adder_IFC;
   method Action      in  (Bit #(32) x, Bit #(32) y);
   method Bit #(32)  out;
endinterface

endpackage
