}�G��J��-�\�P�C���$��+�����̀���h3�ꀟ-+[􈹚���x�i�o�n�+�3G�LF��>�9a�P	~�7��CA�ץ�� ӏ��04u�Ā�N����M��ϡ�^�C*�W=�ho��# ��i�6�eC�R(b_Y���%�X�7��?Z��'���`�J@؇Y�o�L6�~�I@1R��@'A�b�\����T:���~�0��G3�Ρ������p��rTۡ��Z�뤴"!��%�	���\b�	<��,
-��k��q�㳆_}��O�*cTqq�bt-gg��l=�u�M��1n4H�iKD�'La���� b��$jfP��V��k����L�e���[��+֢cR m#���A�q�Y#j�\}b�!/<�Ƚ��ǻ���m�s�Y���˞�	XL�����1�XE���{8u����.�O��i݋��2D�)@�ں�8�OD��_�m�?7�9�A�E�us�#s� |�l�2�G�{��_���8@� ̌˾���̰����xI����g��@�xM��S "�=�V�ǽEșq�f��H9�����,DQ]J�Lw���)�vDO���2��,K�]}��>�5|���ug�#h���dҐ#Ծ}_�}���Q|P����DEXdY�J�^�破N�o#S�4Xʶn���ݽ#�:���Ay�|Te�씲8ENG'{v'���~�-�����T��k����5Y�ޅ��j-R��O D.|2��_˥Q�\D͑��c�Q���"S�Vi�*���)+�;��<Ћ냑U^�!�Dݨ,�O�7W[�Q&��ȸ����ܽ�6w'���=��5Və���Y�_n��VF�.��F����B��%W1�F�A�Z&�5��D\u{5:%ӫ��c8�n���f���b��G�Y���r:�KDe�k���>h�O%P�{k��Ψmj���gPV��N��Z�Y�PBa�M8�!⒟���n�h�F��4�o~�����,a0Ԁnt�
+�c�+���Oe�?5"�����x�]H3���%�ݷ-�6����c1�LS@)�J�O���}:�A�v�4�9��<1ǯ�9Y��Ep�u^���5�mf��`��4��Q�8M݊��Эǖ�Ŋ����� k�Q`�;����<]*�,͉i���Ԥ�|L\�Z��Q�$���nQ(VV���a۩_�����4�h�a��E ��6��(Ce��Srgܜ�+�P��r����=Z/n!�Q����v�A�`�4ɐ�|��I�@֘�> ���}e�d�(��ĩ\�Ulz�T�"��y����u������t�Aʐ�
P[�́xƱzm�k"7���F�Ԍۭ�-���G�ow�۸)�nnp�n~E� sК#9.z]�<�C�"��d�ax��")NU*RS��63�4k�\ޮ�]�K���xq��Ѕ�b�o%m�1��@ރ���7�^�XJ��?��J.��d��f�"�� �6�Xh
ӥ�L`(��l	�q�*k�^������6z����>1&��[�fuq�	Y�w�	-a���gBB"��Ћ�o����F�2�W
�V[2�U6i�}�	�Ȩ��G����Dɇ-h
i[jQ	��:�E��#�L�@,�z�[�a����Um�B0$\��us[ ���u��3�Q����͐�q|A�S`r7��&����z)��6���һ�2#0��{����$Z��֏����V�S���p0��d��G�5Pb�7���i��Ν��~���)}������o���(%FI6Q`�O;��D�;Vt�w[�$�G4��]��iB��Z�8;M0��[˙�Y)��Q�k�^��C��X-87����1BE��1�JҢʸ�]B9j5����ڃ��~���ng���V���ֱᔲQI �&_f�՝���%�壡���E�^��f��^�.���Dh�l�	�5 �G^���d���F���z5�>x]Q||�J>�
*}J5/�U�C��4�d����\����Lh22W`��Q�JK��1c�6i���`����7�o�>���c��ψ�#��;�u����� �{�Q����iф�L�Z(/A�R눍l����,Wv�Y>�^���a�j׮$�j���B&�9��i���Sq3���|�����G��TZE8䙜�1�+F���":��	ѵ�EF��_���z9]�=�����rt �k/m�*ؓ�{��TL݃� ����B���0�`�)k�e	�w 4�HGMC,n`����r=�R|��\2�J���M?�@�Y�=R��}�9�&�R^1�Z���3��	ㆇu��0:���f��Z�\փ��%��W�9��P��m���tW�C}@�]'k�K�S+w+�>;T>>1�u