�VE�+��2��?{	$A�[��6�J�F-�Bgzٛԩ��K����by>pAaTF�]41�낈�4��C
���r$��w��q���Z�@F=꨿��.`���+A.�&�^]�m�� 6)(�>˝Z�%�hj %�Ҍ4�bJ^M|����mϬ4�
��ڨ[�ks�M�Q�q�l6
�N�C��=52w��T�s��3�:2bMZ=�D�����dЕ^!�����-:X��F��h�s@���-���a�m[���k�F�f#��,z��ɯ�z��O2�fY We���{��K�*D�ኒX�ZH�ecdӒ5m�{�5�������V%H��e��5�*o*�T�7��sI7���`�C��ß��=��O�q�sE$��������ZF�Wu�<P��X5xJ�G����ãϧ��s��5�O�c��H�5[�}��4�#�`j�<Y�r�L��cPq��^��_Y���`�c�'������Ǧ)�h	-�����.V[,E�3�!�����H(Ox����bbڛ�O&W�_!0;�@۞�Z��9�.��p^5�F�n���aNĞ�vd�q�Z7����A)�>ҋ�v�5�N�D��pl��M�]R��������?��Z&xj"d2��q���<���YP���f��%o8����Ѐ��f�Q��l1e��ݨ>R�Iv��Ts�21*P�҉�i�f`^�u飉4� ס��+��>H�o2{B�+��6KgN�ш�.f6����‎���#�?�r@e����E�ׯK��ψ����v%���$�L�_�'1b� �y��X�=����ʆ/���eJ�)]1�Q2���s� �)DY��[eA`�,:�[KW
����k����֞%�d��<Vs	(��5:���-Igm��:C-����ŝ����S��$�������/�X�Ά��O�Z ��=�9P�H��p&�-�
���/��&��1s��%� �ĵ���F��'��X	���\:Н9Y��0fр�NS�yĕ]A�T��3���B$5_����D
���jW��pO��H��"c(�O"d�UU^;�����ubn|�	���|�%\	&�d�l�,4�����(�eo+���=�W�@a�hcV6*W�VxD������$Q�@&�G<�`pœ�Ja=E�_H�O��7x�ܸN;[S�z8
��|M rq��Knj�LhO��j�y�*�9�}���'�Ũ� �W-�v�f�u4+�U=?9県5Q� Q��'�5$Ä�_| Zl�=�C��ͺb�Pn�;@@�1��ܨ֛�E�!�(f�H �#C1WGhCz�Q"-ٛ,����H�Ik�ԓʃ��addUt}����D�0"���G�5Iv{�
P�uI��������%���M��q�p8�t��_�E���7e:.#��U 0QCӜ+y*��
 RĹ�ۉ����$i�VH�����2W0�Av<r@���Nȡ-�(z��*C��9��~��j�ӛ��Pn�ܽ�:v���_��Z��8��Y�	cf��f��sY���EW�
>�VL�Z�&��-<�t���d$�1;
L�pAe�BsʫmM�X}���q7Ej�|��Tq��5����c�c�O���N�m��B�gl2���� {�ܠAα�g������e,S����ɮq_�4��r򥢅��s�j1Tc���0�ޞw��h�5@���"��ϘIp�ñm�A�A	M� �9���t����@�sL�2LE�*1��Rs֠[c���?����(�N|l|�AN�.��ޣ��wb���V�I����!	��x���Dj:�:���B������X���B��S����o[̍�U9��pgf�����9�9�e�ZPg�gk1VK��g��7�6�ve��v�G�|2I�Ŋ�v�a�su��W��Va�[��j�)�R��.�����b"4Q��p��S�B懃L�Z빅I��e�ܵ	��P-\a^<џ�ԉuAtb}4�~m��
x! ���]%8��ﳞ����w7�.����D�R�,�	�ȇ?˱��Y��F��$�Ȇp ��BC��}�kNj��l�51�h�@kЛ��Wxs�d��H���Y���l&�둱m�u�ǟ a�g����剣B�b  ��'R��c�L-��������ޘ׏� �9���	�&���@'lp�����Ж�E[}������1�{|<Mr���1*YhԑE�ʅ˪V�A�q)�E��v��F����qi&peG5�>���s!\��Z=F^c�x� H��ظ6�%�̅��Y�	e�I��3��Dڍj��ؕgH��dգ�ۭ���6�[�I� 6�&�X[BWEHl����J�v�3
�x���'�l�笉Jo�'), �(\�^?��Mt�$[Ւ>y0T��]>;�%�|��
"'�M�	Y�^�95���4`�<.�����Z_�(��dp8񸟕&����ɰ:q�-nu`��|�A���6����6�*H�/���43���DE����ݾ��O�Ɂ�`�@�Rd�=S��fƀI��`/�}����s�og�gZ0n~@D���i^@����I$��f�q9?ѿO���)�:��E�Y ���-� �jf�Tj���`/~Krgp�N�$����`5�K53�� ��k� NKأAF�  > ��U�y�<$����@�̻��d�g��0w�r.�d��;�6G3�f*v3�ģCs�ڝ�<�!���Y0Ts홠��	��M�)���`Ȫ��Rm�H�G
1�N���\�fc�A��ėTw߁⃧Dn�Hx}��������4	�~7�
]"A[(rC1r6h���Vu�0�8���e����b�Y��/�׃7|:�k�]��o1NG��%��{��l�i�f��B�k��bK��q莓{&<�M|�� ��lKT考)��$�[WV<��)�P�˫�{W98�L�ޜlgo����A[�9   S ��u�ypN8HPqbD@�̐Ծ�|/	6s[F_�o1ε E������T���?� H�J�stk���On�l"[2��E�l4���k��`�q�Y`��z�@��E�2�4)Txwqe���=��!�{��'��"V sj6��r�nS9%����ڛ��,X�	�{���ipyq��2�x��t޴�j}��h�Y�|kL�wӥ�����j �{��m j�����`ZB��#h��v�+���ׯ�d
b��B睬{c�&��Y�Td'�K��B���1N0�k�Q�Ԑ�P��w�p��@/Ow=(T$��Ӛ��]97ɠVn���#��ĖgyȀ�AH��   @ ��-�����pP��$E2�̞��.��P�9s�nQh9��������+	���o큵�@����i�`P0a6if�i`7Rv9��'l��%�!�7�?��Q2��],x�$搖q���\��-�`��ů��n��*r_�ڜ��o��}fM�Zk�[��o���.�$nM�E�w��*� �3;A'����J ~F���� U��~��/�G�ԝu��U���A��Zm<�_ HK��&�Tî[X���1@N�S�G�����x����*���y�(W�k*�)�oS��B(�uxoAKi���)2���P��z��X�B��g����!��A
�%	�r�Z`-z�s�׫[׫�GIb����T-����[Ƚ��>�D��&!�B@����@ʴ\����Ox2$U7W��p�ǒ�g*S&j�/&�H�k�� '� @��Q�+� |=��@�j��\ؽ���G����%��q�Ǉo���I^�㈈���z���!UP���`L !��Q
#B�X�� |P	� `�t�y�FV"*@g7{8P<�t��霫�f	�d��4A@���U�����S���d[,M��,D�~]�l�
������ȮW��M�$@]{\.mD	��B�{�K� =���si����*wgI����e��R�o53������7�X5ǌn���eE�� `�a�!����D��4E!�XK��bg���i���y���5�)-�`�����/`4Z\]���5���Fs
�0�6�p�Yh]���Ğ�+��YQ[	���`
 �a�
��.� ���+�`�Jx`���+�E�C�x��$T�+�@|X�����V L o��UQZ�q��0 �!���D���<|�0*��e���� `�n���ŝL�����ׯ�!f��2��yvkL�e0�R�ǖRt`F���v_0"��)eI�F""!P�n
(B� BP�]�`�[�Xr�S��־->��m��J��:� ,>�Ӥ�� ���l �| D,���b�B��Dm���ŭl=��Gn��   f�h����C��ޮ��Ls b?!� �F���t�&��P���&\`�� ��h^��z�`lq!깫56V
���Rv��}*��Q]r����h~����my��8l_}iXb)��6����)O�OG�5�t0����W���ڴ���TX�\/�~��'�cj�4v�{�_�T,	���  j&_�qW ���?��/��qd	����Ū�k*�����K���n yY �)��!�F�o6��U�dk��r��3�Q������?���~Bq��^x�_�I!ZB,�l,�񎋪���M�)�H1������g�bѦ��g�5����${�Z�Sř�������v����e�P�����Z��KW�6+��fH� ���KOCI����$��s�}�ߢ����-�7Y��d�y��%\���'*X���>K���M�Ͱ]�L�Ȩ�^�(/�[����OCt*�v�6d�м3�9��}�	�s�q*T%��~���[CH�g�[��=?�5��AA����)��S������5V�l���ɠs^��D�A�.=�����J��=��bg�;n�b���b���]	~D��x������y�g��=3��s�(s�|2*�>��N����a:�^�/NUs�XVrsQ�(	g�W4��=�yk'�
�#�ܬ���q��GIB���R����c�RY�0|�?[�d`}���k�� 