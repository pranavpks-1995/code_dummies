G{Z���7=��>ce��n5�ܰ��[��*U��3ظk<���	�@��u}��Yс`�HQ��>���H{̩�<K�&�3��]?��� <-���A9���UD�f3��d{���L���+�?�epL3>���6CV.{�]%C�D�`i̊�`X��Vx҈M�y�!�.��dcڬP�E�����X������2KeO��	�{�Ss�>jX���4��j�H�D&��υ���x2]:��T�X�@���l2 �i`"�|�R2w�I*�CB�m�4�@ԡQ���^�B�Ŝ�sCF���R���-�\+�w���%EI3���S���������pp� N��FgFҡE.@ڕ����p6���Kq�Ѯ�;L��ꊡ�6�=MOG:�|�����k�9H$#h��g�ǡ`C�ս�!��GC�K�Z�c7����y@n�*���\���7�p���$J5��f[���U@���^M�=~�I�Rrۧ�}�[P�F���@�飮�^X�π|�4�
>��m�?O�@7�A�y�O���B9G�/͙z��U��4�O�?�&q�1H��#�E�6B�Q�o����tF��7�#�jW�Ƅ��+���