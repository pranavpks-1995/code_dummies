package Processing;
	module program (Empty);
	endmodule
endpackage