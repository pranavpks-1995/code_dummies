� X�	d�� ���� ��Ǭ����7���5vЎ<_,���چ�$}���J�P#��
l��F8�G{����Û��.O}�i�EbO�I+nX���ޥ�A��$�by�T�z`k���tx=,VZ�<�7�bw(�C6��Ϛ��wQVϡ��o��#��W��d�$���3�T��:��R�B�cIz�~
��j����J�B�d�"��a�rE�r�22�`!���j��g#=R�����sf�T�Kv��"�=(��|�0A���6^��>)�.v:0���u�K$�i3삖`d�ܧ��E�q��|�2!}�0+*{0@���%l�}U��D	�Ҭg���h�u�Km�͜���x��F���W�S�eC�ekWP�%�e��S��^�Ԣ�ٰ�cyGj1����k&�y7��1��d5��AV�"��$B���pE&�e�'�W���3�Ő�r�M��T@I?��4����d,�2'���3N���o�Q�3�t��.D}�/&lwޙ��}R�MfAVQuӝ�o��"��G]��_C����I��7�U�3��I�D Ȍ�݂nN�>���|���ޜE
T0��.�Mon��i�k�՝�"�)�ON3���
}m�j�$�L�5�9 8վ}KAd�#sr�1Y�a�ܼ(	w��B�$E]	�ُ�4Qw�>�͵�+���) �����/�P�k���5]z�������V�J-N0�rWZ�ش�<{������g�G���u�|OU��u=xm�gg�_9��I��9��S���� �T8��3�ʐ��c���ȁYes�$�pS�u��m[5>_�N��)�qd��N�{;9V1�˗:+U��p����Yq��bo`�FE��n����Y�h�F�ʔJh0��W����/�{h��0X��˔K�k��\�D��x���8J�cLe�
�T�K��g�is.���N��B�1�+�'��N���o�8�_�(�HPoв̞/�AN���+6��F�;���g�UQS[�헤�yL���i���KB�=3��i���8�˂���7���������g��4̅W`m�*�����,�;�d���c��J�f}�Y���T#�F'�"�<�OOy%�Gw%5nA4#~�)|Ҷ���e	�V~J	,��E^�&IC�gO%�TҒ�u�f�u�b�ޙu�����ƦD��¸6�����7�P$��T-T�s��$�k�*�mYUݡu��^Ҟj�=T�u@!H��k60����x*}�x�7�/b�cV�a>�W�F�.�X�g���'�4��6����sR<fb]<U�P���HĚ��Búk�"�8�7��O�d�.ٹz	��Gژ�j�\ʛ^�;�_����SG�K����mr���τ� ��oO�-R�,��Q�������a���7״�<�ܽ����՞������6��t���By�MU�i�pU�.(�j�E]�	�RH�F?G��䱃���D�L���N7xN�_P�t��]��,�a��^��;'᎖���c���%NF�fgaE+����nP�����X꩗���(<���5s�d1OV�o%�T�+P����rX|q�4c��D�h'����QEӖ�t+� �d��4ñbv��(�w�i{8����Rt����yl�ģ��X�0L��LZ� ��)o�^&Lpm �|v�)d��S$Q�յ���q�ǃ�}���st�$��`�X��T���̅~�	g��/,ŒT%Y���ݫ�Q��#�J�&��9�n'��Gt�?A�%)|r�����2���ඤ�P��n=i�}�
H))�;_>b¥�������L�ᖛeN�>���?ьU�env ��{�'�Ϧ�d�lY�#�2LY;��H�/ ��]'�⁵�9��k����C̠���`v�8��T�_�ٰ�
��Z$|�����+��1��5[�	�P?4Kh����?�ͩ�p��g�&��q\3U]��� �f'����W���녊k�0����F)����,��S\�8O����/ɚk;@*$�5P��Q%7��X�8"h������^E�c�)��o��E����?)��f����"͵.��Uk�$�H����"M�)p�cG��?u~KhO�NHm˼��1ūu�ME�8��a��v�C�&E�HV?�a���ox{�y(2 ���Ѐ;)�?ڳa31Boۣ��<������ {�˰s#��p���5�jg3�r���?P�e#�tM�>z����+��ˠ����*��|�Γ/K��df��v��o�P�m��c	��A��)���<�јW�|jIO/9=t�u�	��X9�щ�����э�������VJ�vD��*%��;�Iǒ�Ne��E<�e(��)�@,����u,xP{!��&�y��#b�v����`0ʭ �R���N�L�'���oEK�M�-�>�{����� �:� �͏�q!x��H[�Y�qu��~f?.���?������Kd0q�٭2Oq�k�<�f�_ �Ao�����^��e'�/np4��>��HÝ�V%�9k,�#)DB��l�N2K��������K�f��B���M~P����P�RZ,+I���H7�v�^���P��O�,��n���k���Gh�Ġ��.��\�:�2�G�`V�<�e��ul$�����M��Z����v"F�|-�ӣß�@�g�	���&2*mE;%�QiIj45��~X���Ôs�ۣBЁ8  ��B'R��c�7����I3"

�@т���Y�'�d�7ʌ@�d�RtsFoΟ,������(�MNm�ڿ�����h�����@��0UY�j�~J�n"���%�G�G(��9�S2�0'|R�B�,TW����eLu���3BoD�urMl|�'9o��I��\��(�=#�,�zd� �FX(e�$OI~\�M��/�[�����g��Sͣ�V'H� �c�B,뜕�T�!��w`�at������#  ���TYr�������"݋.1�Zݾ���J:j���X��R����3�+LRń9����P�~�����*:����
��|���siq��^;�'����ij��M���#l���Yhq"�4=v�,�
(��0���V!��KՅvH=���j-�	�R�հ)?[�lO��xJp�����d��M�G0�p�\�s��l��`��P���(�)���|�K�L'�1��}�Zk�����\��H ��%J��������ֈN�<��D/߮�"����%R�99jX7�)Pk/�/���K��o6����
z7��revT}l*�Ӳ(&���/��%DQ�Qr]�F�g��b��&�k�z+��-�E�㠿pSY��c�=�BiV�m�>\�A�ƍ�$k[��]�i��]�m��g�A�oD�*��s�fW�pM�jx���ҫf�d�a/P���]����M��)t���=��̣B4��  , ��U�w��W���%��%�i~��f���4���K��T�Q}�ܙ�18PNc�D��f��8qT?$9ц���/��*ǜ��nQ����6
N请^��4ӮFI7b�c��`.�,�)��Ŷ4))�J����y3]���i��MHڰ�J�DP��g�?@�����ruі1#zv$��{��6�͹;����`7'���t[̰`��ƴ���z�d��]��*��v����[/3� 	�wR�t����Q}� 6"~;��`�.v��N� 19��8볦8�V��`�F\�5�e�h����{�$C�+��YZ:�x|;q��ѷ�M%��J�aȸ��^���rR2C�J��؄�+Cw+���g�#d�>�6NZwz����ҎzZM��/���kU�_A!	?������xe���տ�'�_#�	�]PH3o^�s *�X��A��;��7Z�չߠ%GDM-���  g����Q�p�uП�K�0��`�e��qB�]�D����!
'|��w&��V!��}��������e$���Nk��B��   � �&�u�!���1@�`X.��?���T3�}R?�_Ő[!�a�ȹ���&D���3�����m�XР%%j,��Nb��*��Ӭ��y��D},t���棌f#����'{6�Z��Q�12�?�#w�2R�Q��	�ɉ�L�.���0�Q�o�Ys��9\��-�s�xxIM��!,��eOt!�v1��;aݙ+�~}hZR	�3�g`RY+���'�g���?v��B��gM�K�_��Z��M�3�H�G8�_�9"�#��,q��֣0���u��\8n�57��56����zչIPzY%ZO@�Z�H�Os��B�T}Ui����B<F�mp���'F���9D|4�:rl<�ʅ��3E��U�(��ت~�8�F!X7�5���Upo(�2�� (�z�0 B��^�v�X�����+�(��?�qJ
O��5���/$y����P�����%�+;�N��v���������}��R�U<ʰ�K�����ia���.�c�VWm?�f����u��&��)` �௬;�����#�,&x��̖�5����r%�-�0�sA�l:�ah��CE��3��q�S
R�lEi\�߫Y���;�&�k���n���ʛ��G�u}^sd��0 b���E�<f]����AB�b   : �b-����sa%+�+(HУ���' #A���_,y���BC��5���2����T�JgX��S�����F�;y�1pT�=�4ш���B�̨:�۵�䠧c�cYЁ�{�⋂��#���k���|�gFU�L+�Z����� �=p�^��d�Wr����?5�h���nEdu�L7�G�+�E�mM��(s���l9p���1�L@7�hp��N�oE�L�^�n�F�k`�����Ћ�x�\9�8�<�j\`��X�-�$Gtޝ.���Yp��
���dX�Vr+��6��z����E����������!����!�LD�TP,Lh�� @����g`�K��#�|�>�1P�0�$�E_N����|��S��!�������K>�?:� �Sj~N�'��_�}^6Йn�Lڽ<�KHɛĺ9�Lb���Rص��d=W�]���0�<�Qz�̑�� �^�%٤*�Mĥh�  �!��1��b�H*�`8V��z,���Ѳ��`��gK)��=T`�6���j��	�f��vL n�p��vRO������4`� �^�,脁jR��s�k�ߍ*7B]L	uyV��q����d�EX�.4W-c�`Df���M�WU�C������٭0{��-����h�
�q�k@�٤.����ڠ   �!��0��`�@ p  	H�cƅ�-���"�K�޼s��K	J��z}��U��f���B��  ! q��*� z�,1��>�U�C���r_X�3�Ĝ���!(�׆Į	`C��e��r���� �� @��(�n�wX��OI�v��Gx~�Ԓk��$WT�W~�����1� �     !��HT��7���MP7Z�w^gOC��1v
;y��]L����J4V����7ʭ�-��`ӕG��gx
 ,���=��փ��@*�֎��w�(_��ܪ�b����?���*�   ׍T�n�� �L?];?�A#x�� �I.��x���m�<y��       !��("�%U@(�vk[�|�i�=�^Ǻ/������ц�  ���^���R��8�w���5 ��u�:@���Ք���}K�U�Ut�`������+�b?�tp v�օ�×������%h� \  8��y����� ��>��T��j9��6��N �     !��0��`�@  "�:�)���u1����p\��9�kK�?�6�Z9�xH�n0�	�B0�R�,��Ne� ����{�1Y�������ϋ&�o���%�O����qkX������vx��,�@ 
%��=�5B
�b�.U�L1��	�J*��0    !)��1FB�"JF]h�"Q(3�r�|y�b}p��R�k��B��6 �����myǗ9x�&Kx|�I�L$:IP~(�|�����;;���ֲƾk�i���=A1�o�"#��?,ucB�rf�%ر�����1�( �  K�/�hI)`�@
U�ܖ�dZKU�?}��pv{p!L��D��f���Ut�:��    �!K�I1H:8-2��U؂�����ץ�:r ��1�!�qUg�"䞮Ld�u��7���<��4���k�������V�!F���� �5�IUlbЊ�-�Y{� 8�X�5;1ȗ�w�����u�+2�ڴ��Iդl^����:E&Wl��ȺA�A@��f( �A��@��Ѝ�Z��xH�C=_�VJ��Y�'P����z�{ ��~W����{"��|A+���\USr���pfV�P p�Hρ\   �ֈ����C��+�!���}
e! ����*��.M��pv�!\W2�2#�^�"��~`�����b6�5n�O괊���xiA���H��޾�j��c�׋����(��51��@�D�z��]�?h�NA��O���p,�3�U�U�1>u	s�,@��hj>&Y[ 3�/�Pf�MӦ�cO;��5;��G=%������
��t]N��b�7E� 1;'4�Ys0���b%�U�0p�m���o��@u,Έ*_D�H9?q{�u�\d����!�6͠�h����k�$�o�TlO��ͺ`������]s���o�	ǔ��Dxj�7�Em#P���c���@�Y�n|��L"���ټ��ȃ@~�{����8�~�����P)�)<� 3v$���$v�;w <6e �"��.�.e�����f��,E$��K		�l�X*	e����"�J�����8�7ƨņ7�ٴ��EJlB!�4�44�h���Ji�O!��^��.%���v��X����}��D�����5�}�b�aǣo8?/�`g8��<����Z��M�3�� ���F��T�pDc�F���IL�x-�vǚ��������AR����y� �x|�?(�|ߐ��GF)���#-�M^_�N�K���_�\�%���1XF���d���z&�_��uY��']�	����@���&���!���\Ťk�������T��+�7�/�U
�eR�g�5.��B.lFj��&��ť����)�ؔ`�ἫXV+�e�D��"�u"Rj���V)���?�b�]�tr�؀].;�!��o���+������p�m�ek�݀�ۓL<}�0,#ŗ�:�F`ʍ��S��!�q�p��CR�}]-X�(�]�1�m/�$�g����jnz���&?�i]��1�&&������/!�5"�A7i�%#KB�n�?�\�f)¬��j��N�Ȅ��u!�'�'���}�H&�p�:�)̊�3u>�.t���Ȳ���k�dpv:��r�lc恱�r�d�nU�n�g�ڀIlSvKi=ǜ��w��ӛ���;7<$�$6!aS�
�?N�zqT��U*'����A^yN���-f�t�Q�I��s~�v�����n*0��"�]pC�B9���$�V�g���8�!�~/?�j�:q�Oŏ��l�N��w�ɖ�O�j�E��q��X"�R<%J;R��0�J�N6j�Ϊ6���͐]�U/��C^>禳9��L�*f ��.��m���Xa�7TR؜?sߪ��xj�_����2�p�m-~P���uau���.�^��3x5�2�A��]9��z����۽�~e_O�.k�����	vi�s�R�%�G3�ZjD�NJ{N/N�:������jt�u~<U�FͿ��j���%�;�t0A�YF�R��x��|ӯc��t>��WAQyh:�<;�o�wJ�8��#�K,ۺχ$g6�AU~!���6@��Cw�OQ͕���A[璢��Jѳu&f��4��]%[��6Z\^�Q7��qW�"������V��
O�C�N�F��P����6�����dBuD�@�q|�Um)�<��rf>.�'=��ύ.��<D?��Օl+���7m$͎�'
G�$GՁ���9i�V�ŕ������br�'fb)�S��9'd���;�����$ރ_M�֪(l	�@�&̚�������Ow�C��	{f��2�i� ���!��#�^J^��IH'$��'��-**TA�� @��*4�\��*�;1�`1ۊ�r?�ݵ��j���0_\"��F��$�
�w�ӵBm �nD�Fi�Zhq:.�P���emO�IZ�/Y3+�<�q3�>ۦ��`�uBH�v�Х�ó�a%q�[�:�|�r�љyC��z��F<���Y9^l���h����x�	�����{z@|�;
a����We�+�00M������8���.Q��O�x�s�ni����q���e������2���J����n�1�îjU��k4����֜S@Տ}TJk=�m���x��y[t�u������6,	�����9���b�aN�a�r�(6tv@�݀M��s#����_���~��f���W��={��>��q���;����� H~���5�3g-/ɍ��
��=�74fQ��[ˠѾG���C�$�#p赇i���@4�<*R-*uU���B��	  y��'R��c�3"��P!����@6%��Oڈ��	um�F9Ws5�<xQ� .�Kt�P���K��w$3��'����V�oV�Վ��Jǿ��-���*o0r�(3��V�P�>��?�7/�ԍHU����L��h,��W�j}⏼\��Ҳ�����8��wd�/��v���jˮ=/�o5��]�����\���Ig��i����㣭tG�t����i�'u��5t~��E���dd�P�;
�#�C��m2`p����"�s,23��E��T���Xo0��J�o>��:���b�#��Z���j�C��#P�DS
M��x!n�-�M~Dll��=�^�*�b�~^N���p�Q�
=6�u�!OO����&���11�����F[�ƹGY8�����YD�fNv��p� r-��:�ӓQ���~�.����
"�\��
�L���s��߆gF�C���Փ$s+ ��@�3�����	��{���9��tޑZ��m��.��^B�u=��%0���<��%ޔ^��$T���YU���J��T��^	q¨��z|�<Û��o���z��Z�ث<��ͭ�@����A����=G�R}��Y�����\��A���  � ���U�wn�IaX����;���(_(��&�g�����\�}�u��R���2W�1�m���UC�1	<;�O�"ۋ^vm,4P[��b3+��,�=�;�`�_��m��E�|0L�:$�Ʀ���a�@sh�q��I��{�E8^x���L�\���@��"�l�����& "�@�}h�L����#��;ܾ	B|�+���:����a)�+��>0�$�CPQ�y�Z{V�u:и
�v��T�w4F?�J%�O�'i�&�=휣�S :��3P��i�-��V�i*�r`$s)����̀��Ż�?����V,.�uo81|��E9�ϥ�W	��{�d�w�����G#C�T7:�e:�KE��BG�@��w�a�@������v4�	�}����%e�B@�Aρ�   � ���u�x�ƕW��1�B�K��yVd�,r���)X[@n�{g�l�w#_ �\�{�q50��ܯ����%����9�>���3��8BQ�@��c���V_��K��;7/r�O'��
���� o�������Jྏ� F`.LJҋ���)�|,J,�6)n����pYHWL�aW�B*"�)F���ea�p�
��+B���%7Z�� bЦ��fܰ�>��@�l�����٧L{6�ԥ�s��W�����r˓/^�h,�)S��o]�`D(W@#J��yjF:���z��0z��sp�K�s����.=�kBk�j{�ϣ��q�����!*ְ�J�vy������a�qM��#6_�a3�Cp�R�#�Q�Q�uZ���9D�4���Ӫ�i���? ���e;	���x<��h��`�ɮ����{�,��