�6dZi1����-�����Gԙ.��c�CfZ.����ux�
��@܅(���*{(k��[�[>�5z�|m�nz /�3��1����@�9f�l;�`�	�1��¦m8�H��c�g��F���J��D5_(s�(	霣Fz�  r�'RW�c�J�'�y�$���I����|�Ȳ:}�~�@�Z9�ԞĠ9n��^��'���Z��ye�a��i'cēy�Q��"�ݩ1�i`)��d51��{.��,&�+��O����e"���:!/�T{9�ʎ
&��y3B`�G�ل�sa�[����fP��c��r�^^��J�#�k\j���i�\g��,�^�����Gsf���F]������3��@h'���vw=�x_��$�.`�L���,Y64@[?��R9�V�(�`��#�7��Y"��s�b�r&�N��O?����SCJ�#g� @�B���J�t{��r�#�׻{�G�g=���q���9��UI��R����u	����p�M+By4�@z�^b�k��ɘdX2F	��֦H�2�i��>{|ƟT=j�4�D|��jhHB��5�ѵ�.oBO��7�^��v����5�dN}�J�+8��;п�ff�~0� �-'m.Hc�[�%�}#Z]�dca)h���k�`��MR��f��q �v	����%�������,�;c��+�M���H��&�f,��ILv'ӭ��Ze\����>������Aq�/k^���)��
���l�YS�7,j��a����;�x��r,n���c�7���P���1��b�;�>���D��4zƎ	E�����V�_OJ��o�X�e��d�����-�FF��41G|:جk���옱!MH\��Qݗ��!rw�V/�����YSu���;�T�p� 3�9�� ��(�%���̗o�jz��ņ���ӝ����e`����^""�"���U�lI����d�-�Z1�W��<UTn&��I"�o@) ??y7/��̍���٥�<ٵ)u Df��MR��԰-B�tK�m��F0~��(����W�,?��>n'`>���h��e��H2�6H���QOxdd��r��[����L��U�~�-�r��L�4 ed2�N
˽PJ
-��(��0%:�.��F�sY���͘��L�����Km&��PxL�	�=��{Cb{������g�����Xi��'��W��%���t��Vn8���&=V�Ƭ .�f��5*��(`T�����(��+���c�k�T_,���[���҅��8N0��4����֪��G�K)�.ur5�ۧ��>kF ,YX��;�v� �.BCe B�����WM�f���ZM�aW��,m�i��e�
h�'J#�˫c[�R>�sOM�	�t[���8ڣ���e����t�Ru����O�rc�6�큵��r>3ӳHZqCfg�=@#Ǔ(Cg�趩�{o�2����SN���$��X�[�ѷ�?�/;��zɂ�
�AO��$�%�PH��PA�'	|�ZDj*���P؍5��^��2Y\'i>�z~�j��mOk_���gw4d�MV��;�yv~�8�6
w	Z��Y:FY���T;q�m�Ub�z5p�l�_�-�"���k�'������z���=Y��U��ӣ���eӀe4"�(�ׇ���M*���H*!#	�8ѐ]���B�y)�;������|h��}H�?�k&��G��R����F
�6N>"�Z�Zֻ�Q���M�?�a��W�7;�7 �Cc��  [ ���U�!M��ҁ�dm�徶3������+d&1L���&�	"PD�u),}���]����4\�Q[s^6S(a�>7Ѽ�w��w�p �R`8�p�u��^dɻ�ٳ�`C�d@�8�v����PF�p���X)z�������$�TT>[�"�ihY�1��}f�֫L�o��Sj�UL��e"F�$���\hq��r��b(�6+�(�1��O|@&\.�9�� ��ǈDwfX��ͧ��i�c1j�w�P
�Ǣ��˱���Y��OVʆM���w1�y��Zh��8՞����9h��¢lF�:ʍT�3�<F��2�>+�
Z�$趹�Q���P�]���m9Df����	�G���Q��p�N��eC���i��I��