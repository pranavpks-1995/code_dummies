�=��0�M�Vءpn1��j�[|W7�X@%�)���)7���@�C���   � ��-����A�G,+U������w���"F��	�tN� h�^�G�L�*�N���?�)<U���h��ȩ
��Gv-����ꐗ܅�査��U�98�*�F�`=ܦ����\�A�ˏ
���֌���ώ����&�8�X��-��+���`�Z���뒶���w!���:�S;�FW��ڃ�{B�]�鵺%�K5b`�=��6L ߓL�|����
�pbZ+LC��_��~��|�9��{�&�y����m|��T�J��=��o7ׄ��r}ԉ�p�����<� ���-%/�e%���[v����#V��Ca�p�j����f(h�
遁,_��QHL;#3��L&_"+��y&�R��L�.�*��ճ�j3�d
�[s�I��O�M`��}��(y�g����-���Y�!�4��9$�6߳)��\B)�9U9�3�D�����!ڑ��N�M0橩r]Q׉T@��dOL���dO��C��|��B~���4��%��.��kڼ��*S�d��ҿm-�K?�	�?��L`޴��	�i��|�|Ǌ9(bk,�%�?y�����W �fb	�١�o!*�w;�x:���ӺMPX��?�:9������X!����^_�q��=��j�wY� ыA�w��O��g.J2�� Ε-L��(XWS��"����m
��"����#T���?�2"e����D���B�����XHx%�P=�d�l���p㨽j���"-}D�OQJ=���a�ר3��W�vS�B�fA�sj\�vۜj��4�E�K?��;����!��en<����(S�B_Ö&+q����?�U�([��RӈG[_�$ti��������/���7���L���6y��{T}�+��=���?ˍ҉S]L�^
I�f���^v���УOk��   c֨����C���F�B�l#�������?�6�C_x�I~�E�����F�I�_v����̋���y��HEBm�PĖ<�p��)���M��S&���0��U��4s�����@�0�],�y�1�sG��Ճ-\V�����T �F�͓�g���V�J�y�0������^����S.��f�2nĊ�؀d3���8�I�sb�mp?k�d�8`��\��W��u_���x�19��'yՁB�u�5PO�'�}���N��4{��l�ݲ�:�\���~���f���vEP*����,x�"�d�	�_i�/�fZ+eg�Ķs:�V�0�x����v\[����Ge�S�J�\\�+S+" _D���a�YSo*�:.A�-1�	�b0���%��p��@�/��]S˯�45Cz<���3$��ճ � <fl,ڠ��:������bB�F��ɻ]	�@�`�
�n�@�1)NY^�ݠGe�n�G��c��y�Y�<�(���Ϥ�-V^�ó�+��-�y.�}����)�'�d��&��#��E(� ��xuC����/�W/��!��ԧ���n<E;7t��d8|/0S䜾_�3�����ح�kLDF��t�/��C�i~��hp`����!��{��m��J�z�GB;�.r���H�hs3w3O��s�]�e����|��7��2f��nv^x��Up���#A)��u`J����fYl� ���T�6��� �| h嵘�x?ƙ�*��o��)^�2`:9�1�9o�S��PR�>�U!UlּO�4��I�@V�}�wuz���wBmsjQ�4i��p�_��rV`�u�sf���z9|�I��bBy)��Lf��-'�n�z �-R�U��y�c�\
��0XZQ�h=�ݝ��&�V�8z��^Q�7�dQ9�5�(��9�X �T��b
�V��Ie���"e��,ɝ���E�c.��K)�}Mȴ"a��k�^f�d٥�쵌3��4U`���)_�7� .� _�̕i��Q�Q��H�{�(ȑH<�	�;��FG+�`�~�����FzY�Y�c¿~�}�霅*��Is-ŌC�j���ޟ0��f��%@��,(��kz&��1��ae�@"4�<�󚖌nC3B
Y}��s 졁�-�$�E�cn��W@Z��
�/u,�5���H�j�[��7}��O_f������p�*9�f��C@�?�,�w?<�ŗ��8X��D���O�,h����ē��zqG�άW����m��e9�sV�1�qv�jB�e� :3����	 �~� ~S٬m\� TY�9�] b|�� D���Gi��^oF��Bfj��ܲ`�χ]%S��ߨ�pǮ;b�H^L�u�O{T[Í��4��%c�m�l%������(D!�Ӄ����8�$��G�,��!��HKRy�'"F˂ۢpr�@�{�@�^���ұ4V� �J�;-�6�!�<zu�ǬE���<O�s%��Vh[���?X>�h��h�)�Q���̀z[`���&��G�A;@���؝�T���j�*^]����	�Ё�,��F����޴��T>�^�v����� �p�b	�.���$���ކ{��R��(�0X,�"�JƇ���
��Ɏ�[�Z9�Q[��պ.LjߕRc����JSb ��w��e�E"���[^S�D�!�8������p�V6��Z���%>�n�ǖ�?j֥�Z4����C+")RD*X#r���#�C[���d8�W���/��,���'���o�	��y�]�����Q��Fdl0T���=��e�`�C(��}'O��7z��xOQM��U