���~���� :[X���c9��O�Z��+دe��A��P4�ѫ*D�۰D�m�.5��3������K���X  
"|�����ƭ��}���]�;;�1\)_�&��;!	�HM� rO<�;������4��[��Cn j:�ø&#���qR0�(|�B��Ƕ�[@cK�-`*�BΕ��}����+H�����[���`b#��Eɂ_��������!��5"E� �Yb �p���0Q��&ِ J����[���[�Fq�`@��fa��q�;����ܖ�{C�q/욳ܡRqF���NP�>�-v�K!a�h/�4� w����-5y/4~���Q�E���  : Ej�o�f����$��� Ⱥ��\O9B7,9���k��;&��HAR:+QP !����$�� ��\�"�*8�yx��\mXH�E?��c�͎��������-���O|�Eպ�
LT8ӆ��Ž'�1���a�;�3y$b����2��w��U���y�u_�pcR�L�X Ā  R�hX0�����8Kuyp�i�@?M�gY��n�yk�H |:\T!p V���@*�D  !��9.1��󫫾xX@ BsV��M�F���&�ف/��S�*��I@-@�c[T&��&]�c�=�'ˊ��~8%F�d�B3��F�#,*z��/j�;җ�\1�"��̀ j��I@'	h�Фl�:YMf i���w�)Q0�M4.��ò6�/m�u��n� �٤*�D���� ��!���ޟ���ݵe�\K c� MA�:����"K�t]�������c��x�"����=������/��?&�{p��raB"B5	�f_l�� l$,���8 �!(�|���a]\��X�ǫw�>H��sc�E+J�tϭ�;�i�d|�`3 V�Eo#f����TP�F�!��1"%!�T 
��  %CV�����@���1�I�E��i
>Q. ��:��/|�FsD� ��0��x�g�h�f6�g{]�:��aYH멚��+.��U�eFc$ݚ������M�3� �V F̩���t�Qh_��XsEVC��5i��HR�e�J�ןtQ�� �$M(�k�T��ֈ��  �!��5%#�� X(� ɵk S;Qԍ�-�GqT�B�8��sC�/*���������%�����#B�ƹ/9�Ø��4T`�� N��<�Zs"n�쀤�� H��! A{q@�`�#��Uk�\�:N�Ѐ� N5��TJ�Dw-�����+p�"��i�^���4�T   !��}���:N�(��BA`� Q�$�锈�D������b�u�-gb��|�o�qd�(���Al=*��������,t��}������6�m��2�f�ɭo��Z��!�YZ9 p
]�����Wɸ9=Z��k�NQ��U'����g�y���L���\��t�,�t$ l�T��ƩJ� �!��������z�$ � @%FC()���ht!of�Ɇhk8
-�R�����a֪�C[7*��/�
�H|����ص�,ϙkS�U�#�_\��,ӔKD�x IA� R� S��u�0w���'��z&�� gl�3x��	���%��^�+t��	��s@)K�˖@@^����U�PB �P �a   �0�U��C����
�1�J�nb�*���VRrk�tA�Fw��=`J����L}�^䙐Ye���L~��~8�⬿9�~�]Ƞ��a�+D(��iOûv�n�/�k��{����]��+`c��+�3 Z��\uzp�T�j�� &(���_�ß8·����9�Iu�S��j_ى8�X�,֪�_(�'��޵��؄���������6%' �D�x��c���c��D���2&��W����1	d;M]E/A휪9UN�d����pD)e�d���7�-����M��T��_����P���#�?�5�d꙾�Qf����;�URďռ����ܙKL�j�o=�`���M����d|�Nơ]xC�+�&�y����q�9hfJ��6u�8:F����F��0�hw<Ly"bM<�'��Iׅ�LG��/X����k�̸���$n�sd�O~`k�O��}Ln�C�t��~����6��Dw�_�Z.R��9ϥ����?�9T��:���K�vձ��m�qbqv�C;���<���[�vL�x��@�URpו}j�-z�"���6�9��15#�*��PZ9vf�!�m�_yƻK�@��Q���9
��t|�Q�w���3羐;�g����%��9�t7��B�B�gQQ��m�J�Iu���p��m5
������+a���W[�W��g�,<��0���G-Z���FX�'���L�j�ͪ�#i9�HP�w���nPhE�"c ��D:?䏴�����'5@��u����}!L���S?h�� �
D�"=7�u���"���ML�
���3t�eY�L;���<(����>}˗� �T<,���tM}0�&�)�;6ř�;~�NI&9auX�nՙ�K���@�H��N�ҖHmH����~�8j��b�gHҹ��kQ�j�w�~.i�A�+��7�W��T�1��v���S������7�o#o��ӟk�At�[��ͼB	�ځ���=K�ز�x�6N�$��H�L��X�h��B��c�Ƴ�e�|�����cU!��~y~��ց���KY���I��&H���~����	
���Ϻ[��tˆau	�P���;]�kQ�v��-%3I���u�㕜�vM�mL�7eN���j�v]�9�Oo�b�����qIH1��3`�R���@)�$�ybF١0C\�����MO����h���&x���$��)ᴺ��;G�}�I��C��WJ�*S�l����7� cp��&�^�8P�!�aa���e0*��,�'ϣĤ]4�L9��GT���@£s�B��ֆc������W<c�R�?��.�&�ݱ5n����ɿp�bf7*��K"�a�Ǎ~!�^�M6��*l)�
��^pc}*�c�,�2:I������&k2��-���(�+ �o�.�P�����?VV��͈Y��QC�sƑ�]�����iƙ�xz��EI���uܸ�`W�o������
��(�� �[#�W�&H�&�!��� F�p6�/'FI�YSC��� 7l3���X�iXe��nw�D{�>�v�r�:QK��XR�W���rp���_ ����E:B�)��W����q��f���^o��z�U|
[y��/|9����pI	TS��Y
Ӆui�������õ^R5]]�r�d:Bٯ����Ő(��HGq���uE�"�n�"�;�g�F7Ĝ)E��e�_���kۅ�\,��;�����d�J���꫄"q}���z����?��R�72����՗N�qԞ��D��TG%�����\�k2"��3��lv�������8!A'z�P���C��8T����y��K	8{����$Z�����b�Ϟ����l=5�X�:.n���y/��)m���Y����&�� 1U�'�K�t��?e��o^Z>St����=C/7�i(]6A�_���os�8��t(?����hI�Tڪ^�]��6C�d	����ܜOՃ� Bh��1��k��TQqցP�����Y|�ʂ��
���
	�̓u� k�\�-Y�T�w�2���y2�[XS��N���k��L��0P0cZS��~����+�k�J$ Y
�c�s�M�ŵh�*�g�!�V�hb�I�)	d��-;9υ�#JE�ws	��%�������,��j��4p�ߍx�b`�����	�r��v�F�n��Y��x��fw &���U���ܩDS�Q{q�:�$�?�_�@e�-[Xn9g��a @���!�����hP\D�/������|�M��b^�0W�d����]l���sm��#~H�̥���*�xKʧ��=�kr�k&}>���!�kR /Ā�.)W��J�"�.@�|� j.@� 5r(�o�_(�]s0&�U<o�{��ܗu��������8���6s�-��0u!�v,�h�@�/�8�(�!M	��!w��b��Sʸ�]9Z�R��aW��`�-��6OG�?]"@��������;/#�J���� ��K.����Y�n�s�����|cT�᭄�1?����1��;��(����r�Y�Ӹ��r��=������e����[�i�,�vv~g��mH� ��~�Оۖ�ѵ��Y�i�|K��4���)k��~�ӝޜ2�[T)R��C0�`����,�E_�����
��q|f�'6gw��,k����;��.�n�D��J3�#㎤��r|.��E{�e<TDY�+��$�$��&�ԣ�Q�2�;�Wq����.b�(#�܁6�U��L&����o6��~d�?s<�[�(���`wFuǰ��;��1]�
le<��I��vRO�2 ~Ȉow�45
۱��D������5�p뷐�R-cvY�o�^]�P�����L��>�ޠ;�e{t����p����$~'S�w�� ��DV����Eu��	j��o����k�ܿȎ�9v��|�Rq*r�"�]���W ���T���\��v��1W�E����������b�Ě��|�������I[�Vw��ģӶPzY>X�(�P���98�K�-�p{'�T�W�n��?S��#�C�R\�\<f+�JHN$�/�Hv��Bs�Do:E�"���B]����k[{��к�}Ɩ����ƙ1�]eg��G��D_��QW!;�e��W�*���b��Ra�+T��%������k7C���fSaQ&F�#37;q�yz�����M���J�jkR��-�>�r���D�.��[�N�v
��3�Z�>3��!�m�h��������JM��.(
ݩ�}0�^���a
���M�U�]�� �'C�1㾺'��Ae��12W�l~�Q�R�0\��ž`6��߲�U�VsÚ��m�C���zQ�V����i1cQ�k�fĆ�s�n�Dl��Rס\`��K�����TA�!N7��-XJ�)S�n�Z"�SjS`��O:Q�#G� ���qF�fF��q$����&C�>��z���<]c���y`�y�����6��M�*�;�0����F^=�h���<�d���g�S����B�^B�[�]����=u��/!�!ڿl�L�o7�a��pM�hD*��}���!�H~�"6����8�^��2:	b[5�F���8�{M?*�,�YPR�alL�
˟���I]�����\�0qܒ��j�(�[�{����U���?��w|�6 nK��8�.���p��G�S��L)�w��@�ڑ8�#Q� :"�0Z���,�h�����Rυ�{7=�*�P�ܴJN쮉˩� �UA^��b>v샤n�G)�q��Mٮ�;��>��	���3�T���XL���y��6HEɃ4\}�����E
Z��s�y�QT�09�����e���1ts�w|D.�+@�����A�cKہ��Z�D{��@�1�Bb>z�9��"�7-4<0����~4@3ɴ��FV%�n�v�S�_,`�w>yQ�&t͏ KI��;g�Xݏ��T{�(�����w��"y���I^l'a��D��!c	�¾������m��b��v�a�G�R�lM-
{!E]t����Y\����ihr���`��= bW�
 gAAsS|�w�:[�u:���B<�  4��%R��c�	B����<Q���T��a�����T����'�^�	�M��lQ�N�����G1%F�qw�)H���8�ƈyKZ3��RQg��"&$7�w��-��GQ��>�N�h�8xɦ��T�H:�t�X�D%ȟ9�^s>���򳕕�'E���X�ب��J�����wSY�|,�r	��/-��9�>nX�Y�X���;"�+x��%��-����O"�i(�&���jD%��^�>.��-�U�5�hVbc'��4>�Q:��wUte������:?��Nm�vG9 J�MugDK���e<��ER��Qj����=IQ ���R�F-��$�$ϭ"E��>�aB�Dܶ����A������9���H���4�!4��v��V�Q8�N�a�Ր��X-�_cџ��$A���n�Ӝ���3$�*��(�+�����.b<<��������xh�[���/��4�gi�QƘ=���*F5ʙ=��a����J�؎V��H�Td�_��t��G���+a�3ʮ	�ۚ!����|O�KԀo��NgT�1�������Yܛ@�@ҁ�   � �f���,ta[Y�pi�6@��Eh�5y{��B�#�C�Z��Q����EvM&��Ly@�x(@[\o��܂;]������	 (�bi?%�APAa!�UB�"�U�"EO��p�����C�u����%�i��SS�V��oҀ�����@�:����F��Kԡ��@���Owv򝓦�K�xb���=�����!z��
ʉ�o�ڣ@��7    � ��-W���\a�(��qЗ��n��W��np�kY֕�W���_�� ���+��֟��}�hy@�9�:~iD̫����|���/3f:��I�A}u79^����~���Q}��?��/�ٴ!i`5�J�F��K�㭑�48W��c"ȧ9���+/
�S�-C#ޗ1Z!O	�}}�t|a0@��q9Zڃ~��[i�נ�\q��l����ⷖ]�0���ΰV�g��և �Q��   ��P�UW�C���/��[2E"�i�)���q�4�>���[�:�D�-<7�s�:�9'$ZR��k�x���3C�)��1�q��;�[�����3�D	�P��4�vl�����Ǉ�&7�1���g�Hh� w��1�4��9��H�	`~�l��ѥ=�y�*�VT�Aۥ��
f2y��U�U}��ñNX����Tzu��7���H��S�90���T���l.���=�(����c�Z����~U[�����E1�c�3�����ܛ�ܨJ|���9����@Srf#�ŹoZ�'x4x�ڠ$
k��-��Nwg�e���>�'y���lJ}Z%��d���$�>���>J�r4/��Ik���i8j�]���-{'��0dxq$+B�
0���y��M��ڶ��"���L�}���3���:,��V�;��HG��f�/�* � �)�@��/�-���I��+�a��h��>�<I��{}[�1���%y7T�\g���ò�B@4��^d޺��(Pyz����tn�7�f�:���|_����o;�C����zʭ�Q�JS1(��d^���l�h���4�d�>z�p+n\� 9�%��`tf��ϟܬ�p�<�K*ij����+
�or/�:#RJPɴI�8	,�bL��ׄ�
��ɑT�� ^��- �����z�q+�jv	�����g T��i��|U[�&&��8>\���~4���?���N�p�y�w���v�U��¸�a��l�g*܎zt:,g�����>�^���L����l�͈�~�EyGeK����^?���R+�H �ѝt}Fw5��goޔ]���We��?u����5��R`�u×z�qN�CcGف��#D��6}�F�y������p��T��[!�$�9=�:=UW[t�"�t��(F�o�I얠��X��4���x��l	�n�h8�]���	��_^�u�/$J�SH7�s�u_�Sg�����,��wk\OT���λ�O����s�����^�4��Ƃ�m�������l��
�@�t��E�lQ��r���1QF�,%_�츅�1��!�-I��Ka9�@��۲W�B�9y��{6׭���QNh�����2I%��U,XB-"a0l{��-~���-ֳD�$�z-ⳬ�8i6�X�Jpq;���>	sl�L�1�����iX�yfS��w�����]M�q�P�J��u�f�֥v�X@��Ay��?��#����kR�������vY���'�x���ĺ�zT;/���ݝ䉽4���S��B�ο@6�;>ճ�6+�8�d�T�H.�/��:��K��y���Uդ���#h��l�e���zD����'�ˢi0�$�_��,d��/�Zy%��l,%F���kY�_�B��F�}&v�����$k�	�R��b)=�R��Y����,k��Oe
�'g�V�߅6h��)�I&`�=��p��ua�� g����$��	��e��j�U.�ՙ��:���+�(q�b����n+$&��?���7z�LQ�I>[���cF	++�ΩP�>���R<G?[��g�O���E�]�e�c��TA�REn�����ܧGB�ؙ��b�Bt)�˟B��7���ec�,���+��1"D���j��O@��k\8���1�0@	���Zq�����#bC��w����M��:9:���	�of���������kJw%���P�4�9����ʽ�wkn��BQ_��p6��Xs,e~ݳRz�G�u�(�ՠ�3���5���3�p��"�+�1�V�%_��J�?�3��(C�֎rl��Syc�'���C�0�Z(j�l�g��9�>@0��Q�u䏝ʓ"�#4Wv�QQR����m��Z�yb\��N9?{�	hq/��3U�/E�.�TC�ˣ|,�tlùI�Y�,	�xE�MÆ�蕛t>W�P�+��;�e��w��I�b暿͕r�2��b�=|�
�6kO�\�ڕ�]�`���סM���mG�p�Ր�6�t�2F�"	��U��U��X�_���mp��>��ϊ��b�QP�G3�3��P���lQ�9U��g�\ލ""�葠�$5��݁6z��y���DY�<Tʙ�L��!�̺�
ɴ�i(~�Dp��^����(�\�q�D��rN�0��ߣ����m��)�KH2I�;-�[�!�I��36j�P����5�ʆ���+��R��S<��OlV]��b��а��]��|�#㍌_�ޠD46&�n]R��ۿg-.A���)N��sp��f_�*(��M�Qdsᚔ'vۈ��F��������<����GTMf4a|>f��B���=�7����+p�B��KN�A��\b������42��[���2�K�����8��Dr�ߜo<�<^W)lQ�yl5�����ʌ ��6�NQ��`�~�@�A�na��&E���X�ؔ����	��[��d2ȔG�oǆ��$�k�� ⷒ����5)VT|�2PA��κ�7��{DG�2W���T �A�ӿݱ�:��阞�����{A�=���i0Y��n���� Xr�F���kWr��B��bFԽ�D����������ϓ}sY}xA
�q��T��*��%���p64�n0A��}�i��l���-�U��0b޲�'��ÔS�d���2�GxPoY�!�"1�QZ�vr���l@~�9Bˉ�w�NM���B��k�n�cY1ֽ-bn�^,�"�dO�!��va�.�{�����`���Qi&]���%�ܷ��D�y@����P7���Ѐ���c/(�C�h2?*�l�A�ͧ9%)5a)���~�S	ڡ9>���PÄ��[�#�7	/��c�>�J�q��D@7�$�����y��1�Z�q��;�p7�#���&�+�tY"e-��S�6���Y��ޣ⁘�F��.�W����˰�tA���P��������5��s�S%�j�XD�,�\6Ԧ���Y��l#|Ph7diZ�4j�9ڔ1�Sm�3ť����$�ót�=<�B�+�W�q�4̸)Ao�j�38[0�l���Ȅs��LJъw�d��30��b�i65�(J��1$��rZ`��G��t]X��B���o[ ~.��i& �|�cY�Bw,Lv�Q��}s��c3o�i�9L�p� AM����m��!r���u��� |�TV@x����)���P�����=��b֡��7�Oj�x\��`��#zwz̑]%�� ,ۿK�i����¸���H~oq�~�lx[���}}w�����P�1�%�@:c}O55���>ϑM��h�������Qh�am�7�߫)��tjP������8)®���e��|e�У�5�k���d�CPq-��dL�~���ڔoGC�Xj[;�5�l0`a��`DG���4��]��es��_��l$�q��kaD��)�O��xD������^�|H��E7x�3?qX���T	%�R<$(IM��OM�zP�g@���5��T��֤�+�R]&��Q��O}�+D:�����������I`#��n�NtMR��bd!��y?�����>�&jD����3k��aq��W;e/^%S�[y�3�s��t�PJ��E����������a�(׌�J�Y!ד��S����(1���R%%�;p(�M �ي�k*dܶ>R�A3�bR@SHmjX�ψ�fڬ�ĺ�v[��ݒ�BM*�_�]��+o��{��?#Kg�u�	Za�SY�W�0��	�O��o��6U,���OC�� �怾�P`���)˹����d�oz�dg�9�Hmջ'�����|�J_�/2��°�f^O%�Ƙ�._���!���`��M�}����X/�v�=3�ڳ񧴎-����ŷ��F�:�G�,�!6��Q��6����(��6}�EH �}��4�P�>|b�C�!jq�e��A��p�M�n/�sH�f0c{�+�C�Qg�H![�B��{�Em3�%��0b���":�tc2fG�i�{@X���d��Ih�%1�H�P]�8�(��m���М3��)&��S7ۨ;$r��ԑ`��?Y��̂�n�:�����V�ݓ�@��I����T���U[٨#ʴ�t�ݡ�E=�n�X����[�ɴ�A�lꌰ���ߏ���b��UЋI�	2��{\➡z�N��(����y$�pCՎ��R~�\nBg~�E�Vi��I��[�ǈE�a��S߃l������v��"�G��)J��L�����E"*%�6V�^��٣��ڤ�Ε����V��Ľ`���3{��VbL�S��?��=m;�1`4 �Z��������/ޣ���׽sN���$��c��
)������n������Z�7y~Am@��~�.Dr<����=�w4��7A�����J�/�kp5ja �,����&?�9_������{`�DOCX���B ��  ��%RW�c�YE
`�$e	��Q�+��U�b�U��*o9�I��堝k�;J�<�͂�����I��V6.5#�D����oR: �M+m�r��p���@�y���E�YƸ�`8��i���,?�$����z�~>�E��]�pSH~�<$�S��p�g���[���uBi=�K��'�\�%N��ي%��l@�����O`�����9Q+�Y6�4�8~?���	�b�ʢc�F��F�Q��é}�Cc:+��
wFd��$�b�$�񠻵>�uD@��h.+�(�t�Rc|~nר�4և�3!R�-�ǃjx�#��2�&b�N����@O��E�
D	�����v�i��a(�qC˅Q�m��Uq�"�ο̇/�x�1v�X�uTEMN8w�M8���C�C�j�Z�c�����#�Y�B֬�����Q,=&���,������\�ߧ�,�@|�)��P�8ߝ�ꗰ)O�u�����,�Î���pT�&���9�������@ҁ�   � �����,taWFN1a����j`i����N`!H}�嚕�뚁��k����ne���pG��i<��\-K��.��ˢ����A�D��BU1�f�����$A4�\8�-hXg�~�(�p�P�$� �zK�B#a)1�m��*������ѻ��Q��\s�uH٢R���2�V��l�U`G��Z�H��w�ض,�@���    � �"-W���pi��'���/+{í��{��ٝW��T~�=d���A�Kfo4qz�t��5�y�S��~o�z�8( q�Z�JY�g���򧗧���Y�޳�h�i����`mr�������������<V�$����W����H�@@j�� !8���d��l�
�Ѡ��/v��V�P�n����C���e�}%���rLI
�.��Ӧ�2 ы9p���e��+)�ݤ�ࠣR��   �p�UW�C���0��yŮ����\��+��k��w�z��&�"�kw�G߲���ib`Lu���?�Aw Ҏ��^�@MPƴ#�S��Va�F*��V��4��˷�0>�3��s&�T��b}��4X6��a�/�"�6`����J"����&�0�Ǽ�]2Mf���]X�k�|c�������xCў��V����3κ(�,UC�h�ʂX��9=�X�!{Ŵ�sG�}x�n�u蔹H�;/�v5aY�q]ܾ�|����;��9&�x�>��R��}�&�*'P/�vg�����8��Wn������dM�Í�s������).��@86��\l2!+���A}=���w"�HnZU�U}#���n'/��R���1���-LƩ����ł;=�a�!�_������.b�lF
��&�T����!\�3��Z� ��\f�@�"�O`6e�����e�P@cr@c�:��5���H�'��n#�q1���6
;�A��ߎ#�J�#��ć.��o[z;��3�[���`�ެ��ǓA�r��a�/��\��*�����ʖL��S|z3^l.#��ՙ�3
J{}�̲�-J��v��x��
݅B�N�W�D��Wי����
����cD�@7����̡p��FG�H�L��k��@�l�Y_Dn��&�s�%i=��r3d]P+ʹvb�`�����RhU������X �H��'��F�Wn32�y�z���3Xwe_ζ��?Myݴګ��y���,�E���>�̉uKݺ�E���.�8}��=U�S~�zU�;�ʿ�d�Wi<Wn��u��k$&F��vwz(�7DUEi��'>�����W��|oؖ{���a�|��%Ed$y$
/I����e�Njm���]@��>��F&�������=S��w��f��D?�M5 j9��	da�JNZ�<9ѷ��9W��Ĵ��zㇵvmh��nrA�Z�] xe��M�篺Onްg1��p�!�i��4�)�=L��L����ܒ��4�%u��&/Z�3]4�tJRn�s<�ݶ?�$�2��e��FM��#<�̛��uwTY���q���̈u��<�r�dXw>r�R�9;������,/�D+ﲪ:6k+� 3l*�0S��^���T�ꬃ�q��.5vW�6�j��~y������:1��-��<��>��=^���vi�m�F1�&���a/[���L�Ք��Il�T[ۣwҸd��M���A\o�`wΕ/����j��Șal��%�\W44=�B�6����|�z̀1�ο��w���.rc��
��`�Ns���ƉE���0���G�~�%vO%!��T!�}lؙ�.�m���c�`q.��9�!�g��ߧ9�U�(Ӥ��UQ#c'��K�����-����1��2�;��o"��lv�zx͟�#�0+���E��z]Am�H�џ_����Q��uS�P)e���y:F�1�6H�x�!2��L���4+���R��	�eK�*o�cY\+׭F%+]���q������6���ԋ�SBS>8bXe�Z8o��P�mH���r�0z����{�Z�Yd�Ӄ@�rސR7��@����G�"{����co��A_�۲�ÇeS��}�L�h��g�nL���_o�M�a�,��;Q?y����$39� ���d7�1�s==�}h�.�umc�}D�	ip�ʽGK��j�L�=`�欔)HT������*�\��P"�̫��h����,�Y�x8n`RAs�ʚ!wq�����A�_���N���`h9����=-{�E��:{�j�`)�c�K��
��O�� s�Y�#|�e����^
���[�5�C�\d�(����p,!��g�.Ɗ��}1��^��Q��D�J6@ۋ&�,�݉�r���e�w�Z&��#����Nu)5_���b�v�� �|y�ݛX4�X�k�j� ��rS\py�y�Y(��`	^�����E+����Q�9� �Qk�8Ϋs����f����Nu}�.��W�ty�$h����.��4"e�r;�|��{��Հnȃ6��m�a����$� ���R��w���'�x45���(3IEi�l0�ҙ�\�뷷�;�T�f�Á�@a	�U�=���f���o]�ijjt|/����Ub>����i��/	i���>��
bj�?�H��Jt)����#i�|�W��љ�nc��ϛ7��]<�Q�MTY1r��W dCe�IT_���T`PV}6�8�:�`�3}�x4\ t���QƉ�
���'Ӥ���{;�4鯸����XR�7�"����[|�����J�\&r�5ZC����C�/�a#�Ga;[
�$�Ω��b���V�?�qRS����OYG��-2�*��_�q�]ԯ�u���([��:,��y@r3:���=�}�9���)�]�)`���J_:h'�RJ��]A��^�>x0X�a��0���~����t/w�(D �_E4���U��,֪9�G3���Y��8ޥ�zE2@�|6ƜYؘ:�E��B4�V��Vu��h��+�*F\c��#~�$l?��\� #p�F�}]��b���2D�� ��<E�cD�L�	�Q6�����Q�F#�n��FR���Q��2��c���B�Y�e����/jq��t�n���@f J}���n%�7����e��-s���x�0�Zi�0��������Y���+��L�>�Z�`��t��PD��!�ď�V�]g��j�yV���'��[�Jf�ǅ/�G'e��Q�@�i ��Ό'Y#��
4*�\I�g��Y�<���p߂3��ޞ��T�a:�Β,Wvk�����E�=��@8}\��rr���]��=�I��"��a�dw�H��T��}:���b��$�-���[�ea�Ië���N.wr���<cx-?��������p���&��DJ33�m�S��:(M�M6}��up�ځ$�:ŗ�%���-ŧ�1��E�@�J� ����7��3qt�U��w7n���~�s��]c�1kт����Lx�ȱN�.R*�m��ыd=[\8��j8�����Q���~7r`�:l�T�H�7��/N���������j"I$N�4�*�N�k�i�%�#p�!Z�J���������G���H
�X)[D�P$�Fќ� r�is4l�D� ��*�*�د���U�&[��rzS��Q�3���Y�r�(F��X!��$�
�=3�e�x�e��R#��%�*@w���-��7tK��%���Ὂ�'^;1]����w,��ZQ�_��J�;�&I[ ���.|�#�g�e��E<�_����Wcutf ��=��]zb���D�\ p�d+�t��T{���삣���rt�f��;?v��Pi5ӟp�N���3i�9=w*K�p^p�X���B�"H��S�"FB�Aq�5�d�}���KК`��o��7J�8�^��:�����1,
fy�_nd�"�EC�=J�����5)�H~�fm�ĕ�m��|pߝ�	��;݈�����w]�k2R�'� ݉>�Y������3�k�}��Guo�iy���;[���]!Sė����������KKp�_�nbl`W=�R�
bf+�'	����m�+�K�;��)�� �Ln1�I�B��?�1ىv\t��q�DI�� ��-@��.H�.�x������S0��I�|�=mG��4�x#��GĚDy��"P�c|#L��Uۛ�$$(��"?���P����<��cU��o�R'��7n�&�������Ye�0��(�%���L�%Q�$��2 ��b����a�`�i!s��L�0U
\-�k@����k�~�%��F�|-�ܟ@7�_��;'s�"qj���M��V��#�"�"��2�q d����O
ν7�������%e�/��u"7ގ����u�-�6�w���sI��SIf���Ё�����m-斑�w�GB*�ǸA	/�aڶoI",+�M��=ު�}�Z�U��`�<�I�8�2<�?'����M/�ԧ��j�I`���)�(S�ٓ��RKPmp�#�$�K���࿝�e�̞K��cIFV�7o�ֵ��ʉ��K�� *2��4����%P�~�X$�/l�]�js���<�J˿�K��ŕ��^��fOf5�I`�Us@��\�I�q&^hG�����N�3�:h��?¹�̒��9����9�m���ޛQ`�C��u#S6$T�-���Z,�<�Qk��C׹.���t(�V-��A3{3�W$�ur�$ȡ�T��t������k���fu�u~6%J�k	��l�`�Q�~.��ԜE&b�$ml-1��.T�8=}�Ą��H&��F"������49�h�gN���q��ᖯ
2R����(�dbFv��ƅ���!��rl�G3E�~+*��d����Rb���I&ahc;1���_�N:,P[��W@�� �&��Ny�N�!o�t�۠E�
�����O>	��Y��fl�&[#��R�y�'��}�HM.c��5q��h��y�����L�o��*+)�;�^�Aǁ[  ���%RW�c�Y����*A2��X���yТ��&�na��s4�^���1f�묿p���~����ج����{������v�*�櫑q��Q��a8!����vu�:5V�d�@8"�?P'F�#�V�@s�֩�\Ԕ�P` 0�
HW��bC/�Z�Öw]�@�_Y�W�^R패�t�aZ���Bq���}-"5��*3��osb7� ��D�GK�B�8���J�Eܙ_x�	�ӒF�rv&�P���2��F��᱙.�#�%!0W�|��a���R�I���>��Z�&��+��uCQP��.Q����.KO��>��9��8;
��N�#�#��߀f�ԃ8��$��_n01B�ϴ�������w�RZaIpblմ`.��~���@�u�Ȃ�[޹C,G�&B��۟���4����N�c�o�G�4��6�|����p�@с1   � �f���,taZ��,c����ZU�.KD�%��ֺʎ'٬yA��%,
���+F�wT��t<����$�3P{a"c�N7wzu@b�9����J���t-���m���}��>ܕQ#��/1Þ�A�@����~]d9ɠ��Ƹc�(�8�٣����pz�*;�vM�^��ȯ�T��^��o��� 6�v�3�߭e�@���    � ��-W���@Y��q�2�ĺڮJ� �4��HO9�88�U�׻I� ��Ph3�e�O��:�{�]~mm�lf��|�j�aVH��⅌�i`�n@�L͸�+,-�,�� ,��Nǃ�I�9���sf�w�D�F��5tGzB`fe�ZCTx����+�.PU���q������$B�	�J� *�ʗ*��QR HП�K��}�Ν�p�n�	�J�!.;)C7	����
����E0����������!�������h���pAx	��xok���N�s��Ψ��5H�E���)��\ի��i�Ĳ[$��s!Ա��Y1V�E:��>�����P,S퇍e)��LK�I��a� �#T�"t�L�4OJ5OJ�n�ޝ�r4>ޒ��"F=�2	`�A'IN�	R��K��l ��� �QJ`[����!������- [,�A �M�h^��e�į2ر �Sɤ�ED~Л���M�s�
�e��'�p�����u,h˂K��(O]�盲\�ղ�gx��ͣO@	d9�l @8 ���*��ȼ��`��;n�Y�,AY��Q��B�ɸ@U�٤*�0�J��A0@�!��5r(R�   &]�+����AII�DT�t�Cd�*�)@5���v$0�Œ��0��\�ۊ�i���V�~ξ~����� ���@��&���    , 	Oȴ�`Ӡ�r�i{'�����y�y0�%'����d�{R��f����E�  !��A.)h�A( %�?�[�\�a���-��%��J�	�![kv��S��
T"��len,�zY�YI�,t2VPZ�&���o�4D�I_�'�9/pJ�H�  �,�|���Z3���~b�z70����4Ʃ� fR�
�^�������  !�����&��@�T
�{��u�z�s]�+�y[^/P�2�=��Fu�^�P��u	̬|҅�
�j��� Ũ ��$#v��N@��.T`���"7�fi~�<XL1�����f69�!@  h�A�u!�t��=�HV%􇉙}s�}�ba�K����P�^��I�k�T�Ѝ'��  �!��1/f�
�� , ���W�ԮJ���Q�,S9i��⡈ה�2�"֝b;+�B@����ɦ�С(2��)`L�XR� 4��BӾ�L�iDzE�~S�����J,A
��`�hNiN� �n+J��04�U$Kb�  8!��5k( � X#�2��}T�A$��)��	C#� �Q�
*�.u�`&�/j5^4J�h�����v��9�
A-�̲Se���D�b���fG�ՎI�(SnN�{�I�H�@b0*��� �Jֺ��r����ya�@  �[x�b@%��t�U$0KfE�` 8!��8pn�, yb��X ͟b��4[n1U��Q�+�� �ifZ���{��Թ�6�2��Lޡ ��B�W&$*F��	4p�
#	�@ �X���[!���C���T������'�e�hUY��Dm�Xؾ�tG" �6�!UI	0F��S�U   א�UW�C���<�,E]:*�(u4J4�طdv�
y"�es���@2HKs<������3�V4�(��W��
�s� :Ō׎)�p��J���!m�'�Nͽ�*d��y��.q�'�9��[%X�nGܨ���7jF��'�K�0����FwCuճ��Y�e�
�����GTTA���9A�^�ˍ�2�����qS��(nk��D����>f�Q��.E`T�}�#/�x�0�3~/,~)j!jo'>���[��(}&��z�j�6�S׼
ߎ1�+ZC�9(����5m��v#��%-�q�8�����.!S3e\���!mğh4>KCk�U��O��d���r,��٥��u�g��$�[u�R����;$��:ObYˈ�׃y�ҫ�����+��}#������~n#?����3)Z�jib��^��ˢv0�@�vQG�0тu�ϲ�cu\1��@���p���r#��	:��2CS��9�2BU���"`����ߑk)[9M�mhJ%q� zM!�tԡ){w�71�IYR�M�-�:�Rݕ�0�>��I��D��B�F8��3�Od��y�Btq�J�����g}�0a�l �T�d�_0V$	Og����ܣjq�rB�J.zİ�o�LyY�rc�z�|�36Ĕ�A�C���L��nu��q<�Z?��{�.q98�v�P(6k{�憣{�|�QbK0�E\�F 	>���L��$�qyx�3�E�;9�L�@\�`Wr2r���Ł��ly��F�ܜ�
|���I�g��{��,g�������zU�Q��S����� �Te/�c.$�5i�r0�����[W���5�*8�k���N�P�ƺ�W�^��4 �$���nx\������d*�$թ/�*����*f��{����T��_\By�	�u�� �� x�n䜂�OD����U��\��r�Ca&mCA�$s��#����M�@����Jۄ��L�=��&A���o2���v�_k�bl��Q�6���P�C�֋��3}�O�(��瀵�H�'���L��Gg+�\�W���|cn�_�D¿Qm�C$\�y�Y0KE����K���x����e��"#	C�����vr��\�H��~�E���;�<�H�r�*sL��p ȜI��uO.�Tuc�7��P����ǒJ~pjy�J!Ү�����.��*��t�('6�Wb��gjX5u�( l������el�j��D����+c�8WRs��[x��e���$�'��(\���,��~poT��e6��z0��K�R�HC�y�O����RL�eS��P�r�|�������z=��!�2�����IE��-�>U��yfi�'/�1��V�S{Ł�t˺=����ӆ�"�vP�^�s�����B�ow�mk������[;���,���U]���
f������;+p�IkKj��������FXl~��l�Ó3�s�r�qL�>��M[�=6,	��j\��=ڷ�e�(��,Ȍ�'
?����[8��T��\$�����wFF��G9������ZX5y�J��l���svZu�8��)��A
�.���u����HuO�2���z�$�C5��4��z���]�Wt��d��<]�eu8A(����!�٪���
.�O��y;���쀫y��s��(�clҶ]0�`�aS�]��N�U�#�7�Sv9��H�2ٸT�_m�����*�qAt��p���"j;��Wb������$l�!ǘ�@p�q�?3R���1�]:�!�3�ᤪ�)�[�1����Ʀ/�Q����b4@�0��Q�k)M2x��?Umf�1�3f�A�a$%b���^Y�e6Ӌ�#hj,&��a�$͎�_��W0`���������=K�=��P1�o���O���mz�[f=��~�L�������e���L�c�A�|���nT5��E�w�#m�2�tY��Jc >��}�D��xb�"�Iw�@&�q>�,�٨������M/1�f+m��t	��~oG�dn��j6�E�>{
)���)��� �&!���v^k.�#9��^s�x�a�8%�>���4[^V��::��y�knJ#Q�����C��K�� Y5�H|������[�_9�;8�p���%??f�7d;ۜ�'�a� �,O���[�b��%R[�g�+5�:�׃[���2���Q�^Ȣ�BB�A�!�k�O#�!�,���"ElJ�Cم���A��_`]
Ű�nM$��	�D����U/��G��B����(Tj���쨠L���b����)�8�5���L��T�q�����wh��7W�1֣�z��+�K0z���kL:��2J� \�%��X�˳v�[��{��B"�1��j��I��!}\~�Z������Oxu"G�G;����,��/�ېԌ
7���f�hz-���S��l����U�����Q&Oy!��#Żu��U��_R��;\>ݞ,���z�����XSL���t�C,�3��L�D�G�	�B�XM ⎮��#i�����.�:�,���>f��L%����*[�P0+�>d����y+���|q���\�Ӯ�KgG�M���:_%�R"�oD5ʙ��d4���+fR�D�7�ѴK)F���B]�!���Ъ��#�x�Qf9,�]�Kc������> pLjM>ԽY6Nq_P{AJ.�O�<���@��ؔV�Ղ{��
��|�GR��)B���Gb���c��0�+�N$S�B<v�r����AJ;�ۢjlð'Ή���>��'i��ˉ����cÆ�aK '��Q,�-g�E�z���⒤4{�!74��h�o�J�UK_ǖE
����'}����8�ݤ\	�d�c���iȓ%v�\ת2�7�t��	���+ۨ\�Ee���V����,$�������Bs��5Ĭ����ƴ�c��>:<|9B(y�(�D�<N���Rr��7�8�M�ؽ��`y�;Ũ���/�%�	��\�H��낵$���H����"�3���1a�I]|�M�OM��H��Vg8ĂG���tv��G,�hG�2y(+^�[S�`�r}�y�p[(���-7��]��n���yS���5�1����B�%�����̇�0�z�ͬ~d{���@ܸ��
���0���4'-�z��v�1�����α�l��-���1���p��P9�36��q2%�c=G��ҼZ[xtE.04��>tP9{OR���4+6����

�CjE�vzX���+~�
I8$/$yD�?�^�De�l��a�nqk
J��9q;r���PXb��jt��a9BQs�-F{�T��uILC�[����9��3�:,%�^(���dGS=��m�uaE�o�m�oe����w�b�1��<�	GԚ��hؤs�+�u����ml�B��̀V�����o�.�4�h�x�:�̈^����OZ_� /h@9�k�ͮs�|S���6�fm��Y���3غ~���5Q~q��7��  �P�S|��I��RCSȰ.�%@����>m"N�#RE�p׫G�)8���Pa���'�M�n1�X���,x����,�k�(�^Q��iѱqM/�����--��Y����������,�2�}�OͲ��7�(XmJ��?������`���u+���4T��LB <!SX���;-�CE�_�fb-�"�4�5�G�����yR�	���awO[c��\7���~�"<�O�abwy�p�X���e4Ǚ�v@��,bc�g�.���Ȱ{�0�"��`*��Y(�
7CA�V��R��뎋���[ر���q5���~N���m'*�wV�vBq?Ѳ�X.%��:�������\w�;m��RD�v9�{�4^l`�P���&����?
�iMD�<��`��届ڳ���KO:���z��x�xګ�1�9g�=5�e�c�J���,t����dx���!g�8��]|�<�?���>��D1bL����l@���f��nY�X�=��n� ݏ��pk���S?EF)2�b7��"���_u�X�uK���S����ޓ.bL��Wo����Y�/Z��ژ��Cu"�}����g�����}y����B�y�0De�"��4G��*�Tn�x�}����V����إtĄm�2D��o�r�2�.�V�.�����f8�+h#ٜhY�P	f�	gT�m��x�hB��D:kw�uw��1a�T��?���4"�C�^��K���)^�$�?��4�32=��v�԰���6E7X��ߔ��Dc����O����Bҙ8�V����En�0�t��o!�� �b��"�m|��#�"U�}��d@����'m�=�d��g�m�z���e�,�3���l�E!{�x�3���� �m���ׂ�ʎ:*�	�\���iWs]_�Z����@9}+3h��4UFWy�r�S�g
W���(��~����hnQ�A4 7��4#Zka8�h�^X�R���#A���a��L35���*9�>���	S��sV,�v��
D_U+`��y��Gh¹W
[��c���΍����>>� ��"�9��]��	��@�I8� �B��L�Ȱ��� �
H�F�f;�"D���c@�A�q�p��	����<E/�0B�lU�x��M����;�T��de�V�լm{�f�mA{ʼb���"����~p�q�4�0�ޱ/�O�4�l.@Ϭ�qROa婞@	3��l�Z)'w��������V�j!M����q9L�2H��Fq���"��j�̫2���tg�R��x�����iSL(�V(�Q+����J��УC��  ��%RW�c�G�C3E�"��J/�����|���b���Dy�|�]�	��8�N^L8��U��EA���%9��l��E�Nk*w�Hc6]S���H�n���D�宻���S��x�� �t�7������ϵ�M���\�����a�$*X|!������,�wGr5�l�Qž8V �M�]�=����MoJ����w:V�J�K����&�9��kG.}�t#jV��䮺����V
1\I����PwZ�����j��,���oR2��S��"��lD�`���o�vq���uc�gv4ɷ�{>�Ϙ$���@��6К0s'���붪�Ӏ<����@���d���7
៚�Ck?��/ovhNKz� �2�����,H���a�!ӿKz�k��L�T-�ɋ	�?@����Z|�;ӿ�s��0��Mi�9_�u�SH�� �j2�I����d�r ~��(�`����M�4Z8�7P2�)��m���
�t��)�:��M�wE_R����/w&�n�ڷ����@n�ϫ17��ݖ"�k]���G!m���}\6
����p�jE��A���Dş��ӧ����8�&�=H!���:�4�mo�����]K�^u�+�v&Fj���ȉD��t���@����f��3�?��Mm��rWw�Gj2 Ɛ�	=K�YOP��6��Ke���˓_���s]�ֳY�
dl���3�+�^*_�@�q}*��b�Y�p��-�5���e6������Tk����M4�{H��;j�(��T<\P�/�U"_�њ]-�y["M��=A���~6�s`�@�&8��Q��o8$��>�F���J���,T��/f��e{��;�.���^�Gx&��O�`m�1JA_�ȿU��P.J)QYh�s�\��9hHڳgB��kF=Z����U����F`�q�Aa��  Y �����,ta�XWA5EH��`�RӱǬ,u,R�<��~���s;�Od�bƏ��2�2-���S�7oJ�� `Hu4�% �w�zE�����@���<�L�x���H ��˕`>�7=i�l׍Biy���lHh9a�K��o�8�$�Y���356e�v�b"�B6�VA�$��-�� �@����ܖ�|��5fʎq�lk��w��>n�;2++�:����ͣG��-��Ḱ�:~0�O�V�8�*"�~�)d�͛�򩧏E���dA�kQ_�H���@�9���JHF�Cut�eL&K	~

j��J��:�,�J������A4�jU�� 4��W�� �RNX�4�A��+   � �"-W����B�;D䈌&.�L�;�4J:�+��k���K^=sR��^ú9�>�?r�dy(f���*_�{A�����9+9>�0��uY�a�21��5j�l�����Y	r�����e��y�� ����5pj�HX9���~@M�!�`a���ā~[g���Ӭ�n7�P��ZT&w�)�NF7Hg�" v��W��Hv~�=/�l����.�)�H�n�}D�z_C� ]�c��ɧ����L}>�8�}K}B�t��C6�s���6�Xn�#�[Q�%�b�pS���[^�
H��9	���d���8D
0W\��9b����~��PGJT�Jcf�v̦�z>���e)Ů��*��I�fW���Ń�JEJ�2�S���l��Q�n���/��l@;�'(xk#z��!�aA�)1Z�D�	��������!��0�0lF�(2�M,7M.����Y*|��4]��b��'���0BC�:�g��F��Z��.	�Ve��%$� ��AbC��B@ B,F{����2vK���p���b���<,���L�e�#lT�,.���\��m�5�
�=!DDA�� p!����D�P�j�Qp�_8�7���k�z����3.�C�-r�,����2g,ұ9����e���H^QV0�Ɲ����ȴhk"[=��,
��f��  ],��x{chU����s��K�N �@�o{R�R�w�T�(�d�Z��HUQ�e�A�4 !��T��P�B��k��D��՘0_�"���Z��vXܦc}���wX�Xn��$����*���I�N:K�&S���=$T�f���)P���#��nZ
�C3�����`��%+Ep�@"�ToϹ��{���M�']@�!UH�T  !��-�2 ��aR��` BUysFQ��-�����:?b�k��T�5�K'����ĹN��F�����Bd�Z������-+i�g�@�Zvۺ�q �0��EP XF�u��eh�{���sF`R:;�-pf�H��2���mYX�פ.��Q
�B  �!��91  @���3J
��z�"hy�J��� L�:ѭj�O1*��R�A�OYR9Ij%d�&�BbB'0�ێh�Ί����V�������a�H���]�p
��9h�l�!+��c�$��J�\]9ʴY�v�J٤*�6��0  �!��0t �3���/,��L(��� �ō�������znW�\��Ԛ]f��:����2��T��A	���k�����	#Jd  8 ӟ��d5�3��ȝ��u��h��u�s��ʌ��)��( ��y�s#�H]Rh%T  !��
�<7�  \��W>�5��rǠ��NǶOڡ�Rx�O�^X{#6�����he�W2
'J�(*b�k���RT!�>U��okAb�%QJ$�U�-��{�$)��g]{�-���ϰ�x����JK�&::��@��V4�U)H�[*   8!��<n  ����?`'�u�]s��D���Ю��@
Ν��Y+D���F\�qH $�Cad	N���	nt�Zom�*� H���!B `��mw�TQ��ڝ�~\�~�5�9��ԅ8��"�%xE���	�b���r�K�� �   ���Pԁ&   �׸��W�C����i�M1=,2o,J\�vô��g}�u�VH�f�1�&�9�$9�ϭ��z2~�~<N{S�1O�e\���h92�r2�VN�I�Eb�=�C �|��q�	2C���K�Qh��p��oI��M�+��>���L�YB�gY"*DF�;���ԡ�uP���p���銯 ��L�h�@]3ʵ������;�	 <���}�=P*��U��{�-���M���ȸ9����[��-�ݟP�-�m��7g��t����E0�=��tJ<�/�a3J"��i�j��;S��2^MV�4���V{\^p�=�4odg��UG_|�*Y����O��� ���W�5s�`�ء&Ez'"���Fi�� �<␤fc��s�}��:�f?!�}:��L�D%� �d�ͪB/�9�p�+RМ��)NK��r f#z��m�\�	l/������H�?=._�W@�U��=�+�X��K� v�kx��a%��\��D�KC�	D�4���y��5wq:�yř_bQ
�«��=��:m���|xw�]�	�
N-�.�)���:X"����'�h��9a)�!)7Ȧ&�r^�V��"G�D��j�H��J�c0i+)�v�^h�!o{y�f�A}4-�Ʉ>rH�%�,�*>�C$s�tF��� �e̱
(�n�/�p�bZfx�"^A(e� ^�;P�C!�4;gT�|�,�B�~p�v�������+n�)���t�/R��zD�H9
N��u���3M��Ӑp��RS�(�������G�F�����KG�ܕ�BL�xp����]2D�
-����B�m:��� ��Y/�9�	]�7�K#[ގ@ߠ�( ��B2@�4�e
c�}�a�m0�Է`���W,�K����5�@�νWɒ"�pf
,��5 ���[hu��y�WH�^YUͩ���ٛ�A�A.�=y�����?FS�dgh��2�8�zS�S"1wT���Eu@J+&�����>�甀,ܢ�=�n�\�	�N�|�0D"���?�t�7�j�������2�L���JT�� �	�C|H�'����6c�D��f0ڡ5��'��2s�[�7$3Ԭ8�<�*�d�S�d�ϬU�p�^������D�v��0k4n�SΖ�͇�ı �������/�`����J[���SϠg���E����?.���#����esGe�g��P[���"Hκ��T�h`��0���&;�Ժ*�ݟ������4���ªde��h������j��Ջ��jw��x���k2V>z�����*V�� �;	�/����*r����n�$ +�(�5��iY�.�N�-`�a��S�L��5Ǡ�~��M5pd�h^�N�@���V��6w����ުDL;�'�,��BԵ�;8��%�]��}��3��ǡ\'k9�~�A�#��K}�G]�T����v����OL�݀(F�}s���z6c6a)���00C�@�R1��¡�K����ttV�@dN�9�J��c���u��o�� �%<lW���U�0�!��g�s>����}�R!�o�����K�o��VV�zh9@	-쮕~/1f�v�u�v�+���X�ñ@�7�4�G�E)4����jg 'X����_�����76��V1䇗(k]қ+X�^"m!��=�u�W˧>��pT��^�Tt�U� ���oPsj� �t�B�l �0G���_�ݓ��#C����D���ٰ]Av_�/]�.dY���M:�kP�р9�8�i+N�_�3����L���!�%G�,��K�Օ�� >������l�@3�#��T�)nG�����H��_��P����#�ۋ��wK�0�Dh�]D� ��7
p�E�=|]?�4tW���)\�6�^��T(3�n2e�e��׀���a�*BL��۩,�W3���Nw�����P֘|ŵt�E@�>A����4E�.˟���rW�ϞB �PaI����v�(��>�W�g���������� �'}�(�|6���8S1���U��]�<X��t*35�N-ԥ;��Ɗx��s�$/䞰���S�*"��}���HY g��&P��<��JX�����ܰx��o!��
�B����Ҷ� ;��SјEV�3G�EH��݋j-D��FO�i\cls"�$�H�>��+gι��/+�Y�}v\��� !��t;l�I�Mo��SF����CܲM@X��m��v�"'��J��2�̆�����|E�(�l�6��?:\���:��|	����;0��Ez[	\����n�AD,SMv�"��h�W�%����	����j�ҩ�=Nt��4�q���J��o�f1]�9�l��;w�#]�:*d�l��m�
2������U�fe+�wE��\�
�?���n�	�R3(y!*�Pϓ,R!��ly'�D�oT	��9���SU�(?FoqegUWk�
My1���s4���p�<���fC�E��ZW<�>�c����s��������lQ	�պ��@�q��S�+m�=��#�������a�m������Ui�_[
���:��Mr���B�<���Qr�'�
�\"�[sV>��=un���)�%��0�ع���r�f����V+�z����b�#� ��z_0��B�!�MJ-� �{��<��C[c��f�(�����5���X�A/为�d\���;�D�:p<v[�� ���2Z����q����R�0�÷�eD��Qd�0w�PR���ma�븼�
���-��4pM��zr���Zt㾞�����9h�G_1��:g�D�w��n*9 ɑM�+�}t�𞤟���6Wo�Y���~�k&�&N����Q��4�~&K{���^��1�tZK��[�c�S�q��eMT?^�_������I:�~}�Τp"�袽�}]:�4T
�=} ��Q���:�:4�t2а�><7�RX̋�{Y�����B���'zy�x��9��[j%F����Ko�L����>~M�T�Ձ�1yO�H˕i�=KXm�Z����{F�D�s�Q��8>��6$���W���b2\S�:5-���v�l-,p��$�Lб�\ul�%����P��yٟ����)5en��{j��ԁ��a*j%��Y�n�|9��^����"�mRɢ�:j�7.�;q}rHS�ի�K��w�W�Z+gR�)�����&�J��a�>R2�����v�f|頸+;��/G���v]$���l������e�S������!�M_��j���]u��� \��2�1hhYp���M�ݝ�_��
�F��u�`��
<�����.S�8,}29��;%�Ǹm�/vw�3�j3;��Xԥ�§��X�u��Eu�|�_7H@��ǭ4���u·�Oʩ��}g��[�	��W�͛��8�T1�y𨒡J�������	_�:!�Ï����LvC~��zo���5��U��i�s��B�-�����V;�]�q��G	��j�LoϬ7㙡�)gn$�*��xXd�i�Y��}�UY��U�;��t$x��7��NVx梡�E��e�*��R�S��1����6�3�pA��ΞT�-PVl�x:��+� ���a�i�,g��}��4[Zx���9.����b��V�S�܂yT�Nw�pѨ��7��'��-��C!�<�mXD�|���������!����̆@*�;Y��:u�Y�^[����_,�D�b�LT�Go�j��wP|0�&����V8
"̔����q*�oG{�-mi��:�������-����x�����,�܆�R"Nz�w��0��egbH-DI�j%����Wk�ӏo�Lpj����H��P��y��H<Wz=�[���ZV@�� .����rz$��
2��>]=����]�C/�4u�hb���ݘ�r��^=2�2ۉ�x�a�i#8���G�vt�� ׸X��	K*erגS������-+��������=ha'���[�r��9�Q��Jl�?����MK��ȁ�߆U�z�����OzCH��]`h5/?������:�sY����+}v���r��=��1#�Rj&[�X@uP���0��U'v�A��H��e�sBئ���;Ä^��sS�'2|�[��2'�Zv�E� �k>�CQ����&�ި·'%����SA�Yi�>�L�8�8�T�!�� ��P���`.^�O��A8����B�:��o5�GУC	��  ��'RW�c�e5��3\���C
0�
�TO�8�?c&��4o��юa�j.�X @����3HJ񷲜��I}=I����Z>�d^��'4�{3l���&=��Y���zH��y�0��r����ew2=���"�!�L՚i��d�hÙ�.	)�x�d\ nb6^���u�\D����ž$w��+�K5�E�l��X*�vm�y��$��I����lEK�$��*��I ��eg�PVF��~�: $���ʧ�@T��(\�c�!��eO�;_����F���c~ܣ�$��W���;�+Vz<�l����àt(��,���~����˔��_�ýJx>k��0��$�x��󌟤�S�BA14��J)3���,�4Ƒcy>L�U�LӠ���w?�����2��Q��NI@�����PH�ܪ��
/X0�ײ��R�����$HS�o�f7����s����o�ɴ�~��!&Z�*�ܵ��@�w'�m& �a>B��qk<�$g�$+�g���C�~A5��B7���7���0����te֐_�.�J�^XŒf-Xri����iEh�{�e��=�{����>^�vVR2��+���H�K�?��b�:���:
ir����|�7)��U7+��K�����g��XV�9;���l�(��Gn�T?�@� 7��lPc$�����9[�D���:sNؾC�.�C����bD�D�`Ӌw�+������P(P�i>�+06;���q�����������B�  � �f�U�y(R���ҫ���:�&�Κ���\����~���ak�3�m��fd����Ben�t�dG�z�
�Ղ0�5�^�HF����H=�h����{�IN��.9�����E����i�J�%��q�g���;�z���!���zX6z^q D������4"�ks2��ɧ�H<s�)�P� ����,�4���]#8�7����p�]!����g������l<�|�hZLᆅ��	q?ʱ:�t 5$��H�n,��Rj�	��[!M��1`��'@��#0���غ��e��%�,��!�a5�^�߳����u��ظ��?#�do��1-���n����M�6u���*0!��{S��B ��(�U�� Ч���Z���ǒ�k��67;�6�K�%[�R�5E��x���3�[�����~����[,.�sF�G��M����@�jhkl�@��Qp\��.rp���揵fEwȥ�����f-��[��[���A���   � ���u�w�����9�m�@�#6H�B�2_n�z��ʟ:�CILX3bla?m�1b
˔�	�����ܽ^�Lq�ҹ���w�Yk�g��;$��$vG*�p݆	