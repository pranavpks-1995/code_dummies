>�Y�S*]�;��C�g����J'�K"�2�:�渿uR�̗�G�D_͞�k�LR�4��Cݳ�֏1��/a��Y��`�Z�76�&�����-�ڴ����}|<�t_��@0N2'�5J��֪�A��:��/u,�0���bݽ*��'���$��,�k
�9n����0��gz�D�]9Ħ;�|^9Ŭm+�7.�5(�[��8�B� 2:�fЂ�1kdR�6��'�,�����Ģ�m�,�zy���P�z鏙�����3��	�dh������R_��G��?�FöS1ຸ��
[�/��Z���U�M�9�\�K?�.$�{n8�=�|��<?��M�vtn�ea����Urw_Y�C�	�����P����R��|B,�:�j0�T+���p��ml#ib�����Ĭ
}�n|x�dEI>�� p*��!��
�f_��e��3������l�C���b�	gi{�{d�e,���脖��m~�#� �f7f2��כk�����3����/����J�o!M-q$ea ���mRM�&��rYs����qg�>F��;v�0�S�#��x�g wO"��&��W����2��3���u�}�6���L#����;���:�D�[5P��"�5��!\&靅u���o]-�j�W��ܛ�P�f\���Ȍ6oG�ex�]���%�tEL{�fH�/Kݮ�R	(rѵ�_��{�7#Y��t.��W��|!�U0��ֆ ��Zŗ_�"�zvK@��b��j��p�\�_�"ٽAq��`�Q�W�)�V�>�LWjX�	�����k�����g�$t��D�F[�2.���V�N����������hu�֖'*�-���fW���:�O�a=0cph9g(:!+��EA`3%��1�dz��b�����Ǽ/���Stٺ-�<-nN��Q�(0I�ɏ4=
��4V4*�d�8���N��󥎲�z���E��g�w�_M��2��U��s��؜Ã����G#r$,�&�e^�1+�$=���BT����0+��X<d�"�2�c�0�,��萪���������	�Df��n�N��%;D�����jA$�X��B�Y|Q<ts��amK��S��'@l�QPnp4W����(1�h���Z�r.9��{m0�'l�bz���D�R<�ۮi`^;���̜����M4��Tq;Q<�I���~cZ�8��g�d�`{	Y����;fKY��p��?-�9�Y �7/�딸|AZ�l.%<����~�׌�y��I�.a���}���gz? ���Hz�o�Ҕ� �>Ho�j[�)�y�м��J���y}��W�� $È>�zB�+�Ք�Ҹ��y\2y�����.$ĎR�a%�t�|�/���tx�f�1�T���=>\ �ON�ڈ1����52
|~,h�
T�Ql&�
�H���ts�Ϭ���*�t)��S@��Ì�c:m�gqB
g�[$ �w� Z��!����7�'�(��3ňF'��G�8����m�Z�Z|���$���A�W JÕ;=�� ����3/@��Ȫ*� ō#'� BF�Q4��S/E`*s�K��=��Z�l1��m��Bxސ����BR�����54֨DbR5Sy%ł<��K\X���Mิ��k�����$X�#�Z��;U���۞{�![�,_'�
z���ܞ�g&��g��3R������v	l���n�&��F��Δb�jШ�����dt[�߹�G���wT�Â�n$���b#�"FK���{��hu�oΓa�a��Jv���ߡ1i1͸M	U0�8���Pg���'p�K�öak��aŖ�H`�=�4�%e;{}�I��J/Lx~���&cb�T�Y��V�t n�}g�ɴs�r�j5l�]��-ǝu����6�uܒ�i� е�Q��b��0h=��(�5��!��$4�/AYWL���U�Jo�i�ţ�#�	1#��Ӝ�A=�	�a1����\���أ�f����`zw��Q����ǟ��iE���/7T_3⒌$�.UTʶu9�� ��zM_����$�
0�ҏ}'dZ�R�vt�}wfZq� Px'��Mv��kz~�����n���I�+����x�0�
B�s;{�<�P�5<Վ-�(;��64��D�CT]�6;�0�PZb�*���wE`Z���O����ʬl�=/��;a�Hmj@�F�j`���	�*��6�\y1�/<�������d��Y�%v�;A౱���y�ϣg�#~��P#u�5w����5��l�!D�����߈��>k��u)���{0��|>Z 㡇ү�13��$�f'���aznz}����M`�<:sf�X�v���A�9����K���S�xt&ノ��kZ����;��x��a�b���p�~����;B�iϏcJ���d~ȂE���vFc�w&u�����p���W�{�~������R@�yK���i���+.� ����ِ���l9:����ە֛�b>Gޞ��y�+����	\�9����d�&XO���%�}^��WxSGg�f~�x(ӏ�ૡ�ۚM��זFUU��pXͦ@���LT�K����H�muݚ�����	�ۿtEl��AY�I���D�#��Rp���i�WX��>�7��M���A�cpݹC�oFҘ�&Y/p��p�
̖vpi�|ZĄ�C�b�M
2<�_�Y�J�v�쓡������L/��g4�e[l�<0�����
�/HAε*l��u��S����D\T���[BsOB��?�G�X�Z}c��	V����3APe�k�cԜ�
����D.�$�pQ;r��6��F�1��wxs��D����Ex?��#�Ds㊡�IbZ��s��pj/����x����u�O���J"�~II�u���b�f�N��.2-)�.�6z��nK�1ܳ_�,s�蒢�a]�p�}o���f�����>��]bԌ��g�LO!�1fchN3D�p;������Z��&Ͳ�`e˜8b�J56�ۛ�׾_3) �'���,���%_获(�f5��K3��Y;٤�}��#'���u����c��3��6\9��fy�}R�� �p�{�j����V&7�ʞ�}v�r�Q儹Z��X(�t��6
>9cC4p� ��7a'q�S)��}�VaN����6��y��($�q�E@+�I��Z�t2"�+*��\�-K����FyZ6��S�77�MNU��	',�F ���x[-}Z��r�:G�=��lr	��8y���Q �� YF/O,;!�-U���:H{���"X�Pm
�L�/ݻ +U��˛�����w���A�����!���ӭd���&���F"����;)tB=6���h����o�����D^ ȶ��J�۲
���I�vc��^� G����ot��܇�.Ҽu���$�"��̅�jk4��4X߅��h�|4SO{�x�t'��ε���4^;*�^�*�F�
�Je���	y'�D�@��v�P�%Z�:�IE�������QK�ڳ�{�H|�R��f���[I�@�(�)b�8x���
o�.�O>l�����I����Η�y[�ް���{�%�����?Mv�����dZ��֤?$,I��~�P�giGaW�h���[m�$r��'حA�8�l]� ��M��]ے��Qip���#���c����$�r�S�Z�[4��Y��@k�kԍ�G�kl�Ǯ }d�� -���s���]pU�J������wz��cm.��3�N���