�E��O�	���WY�i)�Oy�3�/�Юn�x�gc���V9�IC�c]r믋֬�*V<��<��6�*@�2�7�r�.@a�7�~�k��_xܐ:c�/��*H�$5� `��qI���ڌa
I-D�!�j��8�S�,�G�4�Mk/�VE�{cV����(���{@���G:4}6+�=^�L��&���Ҏ��������@k��k�Ma���?��9ۊ�j�VZ4�Na����|�.��#�3:4���6�)���)u�r�U��U�T�E�}��� �h�"q���4��ת0
���h��Z�`W��"�y�@Z2lW�R&�&S�.݂M{�Lq��Ŀ?|�^����@��#��{��X��]hM�%@���QĤ�A��+�4���A\��9-��~��z��M�;�6�9Y*�iX��٦u6�̊�x�WL���CN�-����^��
	�cX�E�P2G������[�ט��n�V͠��A}|�/ab���?�L��zL+�IyVa`Sa�ߕ�%�qP;�I��:4e\E� f���l�GB00���ı�����;���s'���_09{���ԃ��;���KQ�*5Y��o����$[�$ތ�7$����9�r�u�J-c��0�zJ��i9���`�]F�l9V��_�(�+#��wOжA�� `��v�,{����Ƃ�/W�p��Xe	�:�0(�=��~�^���4�-�iҞ�)o��ӳ��\ۥ0�
�}������w���S�T��*9��-˄��k�3xn]��G�-�0�����lI�?�- �r��=e�b�n���"	W�Ѵ�ڞ:@��7#�5�D�v��9����皚�f�#����Jږ�ɦ*"p|��� �ydo*b�=�b��� ̔!/�	IOJI��1�kK��Q��nq�����4�
���z�m��:�bv�uP/����\��c�ӥUǽFrR���������V��%Y���nG���o�8��-�ڠ7H����	[P�����c�L�wꄨ�`��B%glzlAg���T�gߊ��>����M��xY�@Km�H��w�E6����Nڃvo��Ѓ��G2|X���i�
<�!'����K�J��`�I�/�8e=��;Gj3�eN�|�G�z:O�;`H�\��ʆ����h;&2\��Q]�9N4���(�.��$�u�}�aJ�F�63�#^v;Wp������~���k~�n�F��!������-}�}^��+��ش

]|����W�R��Ҵ�t>���^`9�.�A��̑�;V��hs)C�����^¦ug�^���a���������&f���G�����^@��ٷ6�qe��_0ݥ��w����ýD���#�� ��U�;"���K�Gx���[�3����s/���(�v�Y��_�����'�]S+���㕓.��t�V�L��N�:M��NL�=,pV�x9x���jr��� zP'�� VWb�z��[�E��4��zl��;�Ŋ�zw[��K�o;&��)KS���o�b�O��2J+��Jzo�ycT�Hn�R-]Ok,�7k�/�r���'{"3�H�
����J��):�)�vH}TdZc��(({���������%$ǣ���c�m��V�$ �w�e715@���HYۧ?�6L����3�Ľ��>=(�n�G�m[�kb.���`�;�f�)���Nm��ڜ�#�*km,����ܔPY�@�*�v�6��OL*�ZSC�-�x�|K�<����
.I�	 ��%��\�3�%N���l��W����'�^%�,&�|�M����%�ʙ����G��;�eܑn|$�+�������[=��wpF���\�Rd�1Wl�Ĥ��h�>s�N­q�[�eg=&�VfϢ"���KX+�-��\��v��3�u3�)�B>TS�Xe���#H�L��/��@�C�c�	��E7nsk����\�AMv�I��R���L�q ��Z�"��o�ָ�;YT�Uk��/�}t�e��BK{<������Uj+(<�j3Y��̒��v�z�
c a)��X�n��J����W���'��8 �.+�5I� Q1V�@Y8H�o���@��'#�ǿ��Cvq�‶�|�yt�3�0dJ���&���/!
;��S��>�m�r�T�Y<�bE��5��]췻"�Ġi���T
-��{��c	�*��>�B0_��K:��[��	�geD�w�D��˘d5�a����)f8-Q�Iu�K=7���`�ʋ��ba{�����+XNa_��f��z%�Hi�,4x���5MH��֤,p1+��ɔ��.ҔTx����O����q�M��P�Dٟ��M=8bE�F1+/
F����.�l�s�E�@����S
\(�d��Q��ڸ�ʨ\��.�;Ic��a�@��=u�� *]�fJ0̀q����CD���^��B���  ��"'R��c�A<(%���������xa����{�|�Z�
�ĜE3���=��}�F���O�Re\_QQ�z��K�w��)�-,��Y/�"�5?����h9I���OC�\����I��2g,�����!&���J#��#��KZ��w`�z��	[�cR��a�s��ד&q��8FV�Y��E�z��}��P\w���>�ȇu_N�lQ���)��4uY��z�&I�Q���#ED6a�Z�����5|�=/��dT�Ej��Yz�j����K��w��=Z9	��:������"+�d�&�x7����G�GH�@������6����~����7�؞�0v@�5<mԂ0�S�w!}-*�C�\X�5n��9jFgKj�8���������혏�z��JB6��w���园��N�#�߀�׹�����(]P4��A�V�ۗ�s�Q[-z���a�Q��ҳKd:Ac4^��a�HZۡ.��o~◳�X��Z{h��-y�J�Q����9��Z�*����u���߈�ݚ�ӆ
;�3[�ֺ���}HԱ^˼�4V�"k��i�2��&|�:e�>o�O��Dp��Å��hJ%�a$sqe%E`y��&���sE����?���0�6��v����d��!� �.�<D�tSכx�����4?��̀		��V�3��;���AW�C  O ���U�uK�����C����r:#Wh���{X�s�=��b8a�@�Nӭ�M���o��!$:O^,�	�����l�j񱀞럹'�r���p��vM���L�v�)�)�95�4��}N� �'��/6�67D.cd&����b�a�h�"���2��K�T-v=)�ٞ������	,'�|�X`cϗ�j��i��X��?�XS2r��Q笸����hE�X�S�RD���~/�����S/����$��3E�>M�xvh��O([�?W�Y�|�A�����ы`�wlJ��m�r����V0v<'���P�P!�Ax�l   p ��u�xJ�"~Ta ����@JeS��pш&���]�\	����*�`ߞ����]>�q�ع���Rp�<������1vlusLuIB!@���k�ɛ��!'�8�K�$'�kB� �d���n�\����Sy����%⒩�ɲ����Rg��w�<ݗ�o����@Gm`�>�G��h�.(����_*C���y=��Eyb���P`
�0�vZ4��?�w�3��ˌ~�?~���Y=��H��FVH��z�D<_�~�(3E�?�E���
m�oob �{��v���#3��x�vJ�Jɱ�e�P��# $�l��n���dH����
;�q,v_ �d3�#�f��F-<�{���ш�`oe�\j�A΁�   � �B-����Λ��!���]R�q0:���Ku����^ٸTDf>?�%���&Ժ�S�l�����~1sI��QĭixxM�	��Dj$���K�uiQ�?L��|�#��үW���g`�����!e?�t�ml����FwO�|����L�̿�n_�֢ԥ�B&�Y��Р�����=?�T(f�P�9c�|�~���H��׮[����n 5�� ���֩�d�+<X`�����1��g\z54��b��M�^M���>ԇA=U��}��&��Y���䱵���v�"�Ԡ���4#<�L��f_W�����f�b9��5��� 5�q���@�{�m�rix+oW���������"�g�M�P7��UÑ{�����Mo94�--i�a�Eު����Ѓ�t��ri7K�����р-��4��[@R����S8�K��@  �R
���`��ER����ĕ���!�����12PY,�Ζ�AG�:��I�>�I�`��,8�5��2M�N���� E7���]�P��R����@�Vr,*�M��+�����EX�ڥ��Ƕ�d4�r�H����c~�{(�cU���{F��l�-V��4��b�o瑲�@K,��P �
 ,4�o���F;t�B���3u��k�&.X� �6i�MA)�
� p!)�ͦHA���
�`,����Rlҷ��Ք\lb��v���p����S�1���^)N l��,���BZ[�>š@	jV�8E{Ѧ�$֌�%�gw�]����G�E�� G2����J��dVhBB� � ,���2ߩ ~���/�����H�g��CY&Aj�a�� x6Pc7~�T������k�!UI�b�J�2 !K�H�b<ل<�h*�p�H������Fh{�.��a[���f�p���$�X}yE%sm�	]�'
|L��X�[��H�����J�ޔ�v;�^ڕG�K��{+���Ij&y]mU_����[�NF����O�B���Zˠ'6��)����]��X���<���(��F�l�T���π�  �!y��#�*��#zS0�b��X����X^��+ch�{���U�
���4�Õ#� ��0)F��L���p]s�9����є���ꔯ�n�����a X)p&�A�x���)�UU+Yq(o��|�(��(^��Υ=x�  !��Vf � =�z�%��!fLhvߵ�A�8t:cg�s�#w�u�:(��l���S�����3��1��t'p1:�r���Y].�6_|I~��ҹmH2/�oR*��Eb�#�DN�>0���
'j�g���P���n�,�[�/� !��T� @<�U�f� �����K	������ɭ���p�j�/w�de����_�}�쓏F���ܕ�
v;�����3������m�h=�S|-v}��FՈ:���+��"Ŧx��[���"� A-��t�+?2����� 8!��X# �і3���]��AR/��j�`3����&�:�w�pC�Ó��������oO2Ǖ�;��2+@�c�"����1]TH�C)��]�~��^ٯ���*Lu��p^(5�|�|�Cp40��@��I��m4e=�HUR�ܱ-�� !���Ff��L�,���5�Q��lh��.�'6I�6�󘟵蕿�A��k��i+�i���zm�q�I�G��'��$9;�s���_(���jH�a\���`k��I/֧���- 3�D��K�� ��� 5�B)w
�"��B���%��QG@�M���   �������C���U+z�/E�<C�����;k;�9nn�u�-�e�S���cu�2����g��)�{�2�Ǆ��M~����Q;̸"��ڵ��`������W*ς���b��M$�	�5!��j���m��~�#��Rc��fl�;�r��d�n���c���r*54�ā�硡lِ:O��e���{˚4���B�
d�'�0z�j�J�d?F�6�d-�E��Ĝ��C��䝴S��t�=��i���5��p(���FK�`hN*�ɤ&	'��^�\}�5Py�fAY�X![Ci/*���*^�[�Ϥ�=H�Y�����Bz�^	�O(�E�أ1�63��"~�j��9IHJo3?�|��>ڽ�(�F�`E� m�1�'P��Y]8�����Ӛ�&��coK����Zv��u�7pS�d4�@�����i��iP�IV�yi̭FEd",?g����`ȷ���OvA#��'�����|`���q�A�8qO��ǯA�,_BE���;:⯆h�]����`F\��� ����QQ�$k�e���ކ�'C>�&�=����@�m� ����ԁ�M�=T켱�1�IoNV�����������9��l��.�l��Q���^v$�V�G(/��*����%Zĕ��Lw�R7�R
/ ap���؛ ��T�%<�qP5�Ď�P�e���^}-�,-�H��m��d��
3�@����>Ă/�����H4�#�	�p�
5Y��b๑�-+V8;�i0���x�3�@dl��f�¼/Nք���]�#�/h��8r��b�CB�;�]��Ü�y6�p_�'|��a>��	y%Z�,��k��dR������J	H�0���܂�X�/nO";�D$�1���m
=��t��Q̒����������d4;�P��8����d�'�%MH�h� �O��ɺ�9hP�����A5��Pu�5A�L �$t��#��;Cl���,����k	�m�������hΪM���y��m5+}*)O�P���<p*����iK��O	(L>h��׉�������>�+9��3���o�@���\�c8��CMy:0���1�sk�fe�U�/���ݡ흄6ܯ%���6����HP������gc������~�\��:�D#Nٛ'�$�s��ѝ�b޵�m�����+�
�)�����vX
�V`�����[�]����\�%���q6��#[��@�N�Ύ4��P�A�^�d����i4E���+�#����)��(�m=�	HC���dm'�t��D��o����D�C
^d@�����8�Y*	�閘��KxHy���{��ѓ�0�Ғ�����?����s