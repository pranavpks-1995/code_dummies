iC�%�o1� w����aJ$�v��m��a�
\�(�g`�Ҏ���15�i�c�{a>'�E�����w�0���o�~�
G�Z3f�^	[�lֳ�w�$)��Y����$|�k�f�A3���y��E��/[�A+x��m�}F Wkh'qsC"��q����P�ڢ�7OL��R'%�v~�<Co��yޥ� �Ncc܇y�{�~�&4�j}��r�W��=�}x:��K~�}����>�$O���f;隫`����۔�n��O��Z��o�W�?k��sl�,�^�^SF)Ū$b|Q�n>�
&�+���v\������Z�sl3�)	oԭ�'Se�B�!�B�1�+.�fNA�^&1(�)�|Ze����i�8�| $ �t�2��c�ՊV�V���Y��;<������u�g^F�EzgU��4���@��1�!����C��l1�[�e�� ���J%f.�_�C=U��ݺ�)w������߅o?�u*�v�+>�F��+�Qv�{�����h�A.�7 �[h�]B��ތ1пYY��U�02��+F���@ �}���@HG
NJRܹ� &�AĦ�,�j���.٤*���q�`  �C�u!r���� I��  �  I�*��]"q�����=�mmŵ�UG����C_D���t�8��-t(Q�ϔ }4��_a$��CT�xAq���-i�c�D�9��J�)���_B�^�8�E[�r���t�'�q?�}�u6R TՏY�����G�d"�٭�}uh-�@�����q� d����뇔�A�bu�򱖯|&o�J͋=u�ӨPg��I-� cAJ(���2��C��		G�P�N�VB�g��91z&K�r�4H��)�_M߁s�Aӣ��]��h^ħ)���y�r�R(��-�j9�J�y|���!F�r]����!���h��p+�_�k.~e��G��&y�up�H0H
G�g�X�E�=`@�j�����~hNhPr��)>a���3�lZ��Y�{t�'���8�2xt �-t�X���5
� T��E�#�;ӷ�~�ʥ�Ѧ��r��P�\�OE�x���,���d:�Vܚ�-�Ń������D��d��Xcz�V,1ݙ�1flN�6�0�8.�ɐ�/�SN{�M0g��\d�О<��	).�����2uA�5��ȼ�?�A��&f���v�K�^�1c�oim�WJ�!��,܊kc$/(̡��9���,��)�w�k�	��I��2Wp!Y]�W�c�ˍͧ���C�E���
���d�����zO�
����JKaHO������X}�d���3�x��r��#6�B�D?��^8�t��&1T{G����E�k��v�K�n�,V�.�47�ɅH��OrQ��hG���}��f�Yܦ���|����2rѸ���������'�#ހ�h�H�aŮ�"�o<y7̰�	�D���E-���z�I�ҵ �f?KE4�)�z,�X��. =۫��OS!�1���;�	Z��qb���cP��Y����GZ����L�=�v�IJ���A
�(��?ΧLN�#��r����2k�7ꔇ,� Y}g�\��H�<�BE���˹Ya�^�!t$)�P$]f�-������#�4%�k�Y�"���##x��y�GTŧa��p(�m���)n�)2-;y ��VJ�4�� C������o�.��r�J��:&J���=���N��_�8�|�d��[�f�-��u;'W�q�ۈ������`%׵ሣ9~