�ҝ�Y�;v����<�_�q�F�O�ߍOB5�aO@I���u�b�0ߔeV[������SQ��*<l��t?��~�j�z�H������M�(|`ЕX��4�moZ2��؃�Qx�=.����X�\�Gԅ���K�y>\,�,�o������U��"�d���q]Ek!��E����<�\��טD.-,�1�gE�aV�\�ݎ�9��mq}"&�m��)�m���	�V�«��:Y��������0K�6�hY��|�c@�ӳ�?@NX��@��{���Z2yu�BxM�Ԗ��#i=`;���"����X�)�%���^�?썤�٬o-�Ur�x���0���*X�8�Z@a�᠞�B��)��e}$Ŀ�,{v9��vAG]�{��2��ζ��Kt�� ��K�����q�����ֿ�ִ�vW�l䒺�� �X�8����(	"������>���1���}ئy��JkF�H6S���S����VY_�|=e�0*u.,�N��������f��7�r�
�� ɾ[�\��\x
R�ɉ��іG����V+^�0����"��;�94=Ǌ-W���λ3Zq��<��/������`1mV���_�?�9Y�"V����H��=,-�~�	���/4��ѩ�:��g�cZ1���7�L