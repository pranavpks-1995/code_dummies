��9D,�0��y�TH�k�~���0"xf@%�"��}J�'� ��}�~>�~�>�&q��/��pO��c��+�gS�Ή��#��Z�B��xv�c������_�cp�񁪋��w}��s�� ��-�+�����D��p�b�/�����H��֮U"�\}3�k�;4a�lq�x��>�K�J��h`Vx�=6��H���;黠>Y�G*�V'���1z�G��il�)�ϓ���$_��O���3��wz��<��&�s ��c�dG���!3|
�}�$�|��Ks��*3��3
���k��sF�!(�ܼy֛��\���x�OqP|Z�5�U��A�CV��u%Kl?��R��/@�d,V��-�t���}.S񉇺rB��*�ݬ�y3�t�q�lp�����R����t�VE�o�����=�'�sA.��F��P�Y����(�~�߾G�n�d��O!�s/׌�C�c��3I�� ��A��ag���M�G])o�|k'Wd��k�_q��J��)j!��d~dw|���d9'��75*��suaY����m.����ȞQk٣�O�}.���	ٸ�>��3��!IҀ]#�*�@��X|�r�mR;7�j��uY�QX�����϶-m6� �>�r��{wV�Οlw�S�e'ml�{����?�i�ħI��l��vP#��/Rݽ
�2�O�͔z0��H!W�U���mU����0B��"�y&]Nd�ס8 b���6S���j?'c���Ku@)+��/�pM/�W�;�5�c,��g\�9�i����Ig	W!�R�>�����Pp$g�)��� YH�?!�B'YB���)�,�Y_Q�!�i��4!�.f�g�	����R <���4�T\\ÿ0��8_��t	n��R�
�O��P��|��/6uH,�O������a�}LU����;���]&^�ɚ�G�������t����2�V����d��\DnaB<�I���r��I�:�²G�V!��)��c|X��$X�����V�*�q��[��ۀ�?h˽%S2��SnI7ǐ�ԑ���^���jUA*\f��� ���}������	����p-\��MSH�	�h�M�*���g��y�p�.)%�5#2G��[j�R�Hʌ������Lmy���:\xUEOs}��ތ72��,�e�9���d�n�#� �nu�=���Rjl�f��ɐ����4C�s3��C�\��7�Dy�C"�� ��+�w�SSÈ���dN���/��1��U�ր��r�I/�Fx��j��~�"�\k�4�X5=�f���`{�-���^���NBCA��8��K$��2�v����\��Ծ�>��/�ϵ_܄�^�Q�� ���Q=ZP�hE$�Oݠ|�����4`4���E���'�G��@�0x����߯��)��=X��0�XML:��`,EҠ^��
����@��\a%�mY�$���;�^_�R�0�%Q��=��9�����g7�&�O^NS���q^�p���m����ƃ�"hM7��"����.�ުb+~��]}Hc��z���p�J�b�Q���S�֝�ޥ�L 2����A.�tbl�u�p�E���r�.�R��Y�^!$W��k�*��p�1�;mD����P8�fG�T	�h�gI�E�V�y�yO�"�5H��h��{�q��� G��8 V��Wa������U�г��j�
ճ�YU�̋1h�*="m�%W|�;�(@#<ޭ�#�T6#AԪ��w�B
��,��]t�F�)uU|�Z��N��9����<V�rN�k|[W���Ƥ�ݝ/6Q����I��84����^�)̏l$J��������I��bgs�s+ۭ���!h�����p�\�`�7�XX#q�T	�GQ��MGQ۞�0F#&P��;��!�C��Pd7�Ȓ��l�$Qp!Y=���}�v�G ,- ybJ��߈�A&O�@m

�.���KK}����W+V�
z(��!�*هvo얎Ih�PLL��P�M_�q��D7�.Bt���2�	�`T!^��s�|3��VQQ��I��m9�P0U�',U'n�.�I˕O;�{L$f����&�4�˨åJ��3��.]���ҭ`��/��^�a��%ڞC�V�0��(T���cֆ�[G�Ջ���!`��L;b��v�_�m�*?yX.�ւ�-W@����Q��я�2�3Z=Ps��$����2���/Ϝ~V�Z��q�/��i�2{A��}���v)���l�v?ܮ�Ċ�c���RZ�r�90ܴ�؄"ԭb*n�E���'�|8(������_��3g~�Z�r.�h�z�4����.���� T�y�EE���8�G��cz�+&�:�%C�S�\c�#��YA���=�ʓ ��Go-@�x�$����}���d�Z�&�ܔ���$����>��܉y.�1�6�ؖ���PI��B��[���V���V'U�"ut�1ui�+��0�%��;z����<���<��9ε����뻙�L6J��,A�G4ċA=�������Onz�; DJج�r�`�c�r�'�=툕X��hi�֌S������+�=U�׵CQ�T{��l����<����А,�d�/Uk4=3�����������&�m9�Y�PxJ���R��/���a�1v���)xh���J2���omA�Y\�f?��pZʻ#�k;�Aʙ������D�b�Nz�U¼6�hP/{�6m4�2	���ӕn���`*M?��11�_3�Y����ѿd�p2
�Ϟ]���v.�av+6U�0�XȪFl����'�Y>��8#x�ry�Hk��O$�g�d�Ѓ^�:�X������"����p���ӒL��:�2�� TD?��*T;!�*�k:FEv�+�<�����l�7ûR�-\�b	|!�^n بs	愬3_Y�Q����'��{�,�����"s���u_e�l���*}���\?�]u���M�X�6�T���Z�Ù��h�T"�����AKnդ+�iB.�����K��u��v:��K��5X^��V�"pd�~����+�Cuv޶��  =�'`�Ҷ�`ơ�>h���H͏J������<�:�~���}34&BB�bh�����>��!Σ��rB����z��E.vZ<`�-%{�1�B\q!��Ѿ�@�njn�C�����CO���,n���~����nm�~�����h��Mӣ٤Յ3�H���%��e{��ۄ$���<
YXI}��4����q+�1zWݤ�gp�B�.NNĠ?�Jᄉ �I�(�t�A���D�Y,�E@� !��������!��`�s��
�T �:s���Mk`+�
�Z_N�jX"ѧ���b�κ���[��PL������R|�rDX^������RD�8ll  X,B
̾���U�}j#�&X��"U��ӂ����C��+��|s�yE��)�P'R�-q�K��T�3(�p
  �!��!��Ȉ!�m�h`�C���Ќ��z5�LV����XD>��Y~�����ԺW���IXGI4�Yi.u3�zr��W5��u�K ��-F�`� 0�~x$5�@�Y�����"�È�ji=q�1M�v����pl�Q)`���vJ�b�P��HUR��T���e !��w��l�X� j��І<{h<�H�mjH �b��f�W��6���U�����/<{֋,�XGm�gDfB��n% ?��S�?Y&�#X�(�` , ëА��QW=�C�qAd�L?C��1��[��J��^Ⲯ�8乯j�V�l F�!UK�\���� !��0X �� �E�Le+h���7�ڡ�������KPMX�+� 	�� �@�JQX�P���5  ���-R��)>���s��	�/Ć���ӭ�1'�D��tչ&cae������B�_Z�����A 	���D�m�T�"й(1��� �!��8Є  �
�Pu 	�q���G�NK�"by ��Pf7'za����J������>���Z�k� ���!�>	��b�O$�Ad��XN=�� 	f"0X�	�  �����^L�|��0~��'y���.熫�c��ӟ@2&�"e�n�}E��Vȗ�oM�K�jÉ�m�HURʅlj�	�!��0�3 e�e/EJ,]H�/��GH"Ri�rH.�^kѕ9�䩺�w��9b�:�,�r$��cu���FA1LJ^Ap3	VY�) ���������d{q�d_�]/7�X�9�,.��C���Pt��� �d�%6oϙ�a�z�o�^���VT�(�!��
��@�/&�dEvƈ@j;4���u8��\Om����I��JF���U<�gJ��hY�96l�c�1j�)6�ގ\/y�!����UM�� �V;<<?V�|������҆���wuz�V��^� v��1�M{��� ^ �:��@m�T��4� �!���B�@�Da��p�W�޵*�(�hѠL�T<g��?���7���a���3g���7<3И��~f'���J!U��7��[�3nڱ>ZR5A-�e��],80]�@�**Z(��F���\�MX}DU߷HURhw�E@a[Z��F� �   ��I�c������D�����(-���0�g�P xIP
�a4,��̂�غ���I%�E@�e����t�Cf0��`p����k^dC�>�R��Q�~&sw�no�C���Y��W���h�]��;6��֜펋��tW��xJ�G<l��im��*9$Շa����LE��~��ѩ|i����@�^�W�]I���|�Ln�{l��*>��u\>��1�Y�O�����]qa
F��O��E־���)^��ٷ#`.#�?C�{l�y�`�vJ3��~xà�F�:�mŰ�+��rT��	�G�v����w?pf��bnΠ?I�n��	?�)*Ƴ��!?�8b���C"2]�)��� ��\e*m�Vq`>O��>���C�P�
��ɣ��D�o ��!�v��j�߲Xh�c�1��Ь�~���9�,YC��J�(�4R]��}�sO'��T'Ӌ[�j�Vo-cI]���Ax�Q��:iG��X�;�\�E�Dg`�~�k���kH9LV�9�^�+�N�J���+p��@���w�aP���gQ�C�hiD���0����.ݭ'����*)�(�t�ù�,���4^�W�0(���l��G�ah��0�Js��1�(1��c�W�u+=��æy��P��'D�߮�]w�D����{��&��1��$7��$�Xc�>w��*�O��C�3n�W��P��\
L��*��_�����恖¨�ox�A�W�ϳ�qLY���:xEְ�+�`��_��y�M�`��f��
�˳L˅`��`�����ȝ�ԫ1��O g<���ϔʔ�dk}4�^�β����}�U��Ʉ�趹�^r/�W���i��c3�A dg�&9���
w:(Qyy7I���\�1��;�����7Aĭ�ZЂKQf�.�%�桻�{�@
J��rУNf�KX�_���څt|X����X^�9P8�ÍJ�:�3�oފ�,U2 ��"W�ܬ�m�^����\t k��T
��zg�4�����A�N�#	�e�]��؋w��5"W���Z~o��y����ۗEO�����`��m���������g3�X��~�>ϙ��+��L�#;���\��KP���Ж��%��Z��8��Pe�X�R3���h,�,�rX�=���[(�
��ʋ�@H�Y��H���{���=<�����`�O�y�r�/ۨ�V����}L�#PB��R`n�1F=��g˻�uҾ��ݻ��kt�M�\�g`{s���o�$X�d��z��B'ͼw�F�^T����ߨ��J���h)ıl�V7�"�#©��ddm��Y�q��l~�ev�t|\G����Y�!�L
_�^�ے�7J[3Uc�V�!Bf��� �瞦�%p��S����i�f'�����n`H�THHJ2�p������\���-��֧�N��������I����h�"!�9���!���<�Ӛ=07�J��/a�����#2�\���F�_��,7���]�Q������Gz���h� Xj�5=����
��s|>M3I$�Og>�3S�����H0��f�/ qe$��^7�;��S;dV��%%�<����aX�K�0��X�'�Ⲭx�%E�e(�ӥ�#G�Ed���R�e� ǭ�&6:�ל$>iRxR���C#��y��@-����b�x��Eo������.�M��,0��ʥ��wƔ��n%��NWq~y�4�j���s�LA����k��}hz�����N���n�A@� S  8��xc�p�e�4,8h���)=R'��!���H�A�~�n�H�/��nxk��M�[~Y����L"$V�e��R. {��@�N ��E@"���8Xhn
�Yvi[����A6^�r���e�KW�ޙVyb(KB�,Ud��*������fD�vZ
?���r�4�Kt=�~���3E<q�V���/$݌W�XB������(9���>���O&Oi��eګx!^��� �5���"6�.G,��!�i��y�5�O������U4'X�P��]��`�@-8�F ���߱����nF�����Q�����@� )   � ���~�o& rJ1�&�a����Ȃח�#�h���qp{�n�a?�H<[e�6�v�ZLjWIVo���'HZn�!Я�{g:��g�ڙZ,d
*�"�a?��#�#�m?ɔ^"��h��3��7�,�B+��pG��d�E�S(yO���"��E�`�dL�W&03*�>2���G��v��Xe9DZ���a�t �bEq�}��s@��w�[h� k~G���6P�A(� }     �&��F:0��fT������$��oq�/��l[�_Z� �R���|���!�}�#���R���b2�3 �m�6&��0�D�t�O��>e�	6]]�h�b��4/����
n>DJ OQU��*�n�%���I�$ կ!k{�$J�y��/jYՃ9&��Z3O��kBt��f�6�ZK��� �˯.�~mAϨE��Yn/@!1k;��{@�ա��׎@�9����Ԁ�X�"��[�r��`&�@Q��/ԴR��~^��H�k�39� �C�.�e������EH�v��������!������ R��a04�
��#H�O/,���Ru�<xa�ʧ��/��ڮr8�2����z���Y��ov�k���g���;�N������R��8?L���N��j��^�$R��^ץ�˳\����ڠ��A�0��[i��U�����r�4���!UJ��l� [;� !�`FB AUVx ]�X8�`�^w�@
v�=��y$����n�{;3������I�q�19����u�.��g�3B�B��柇�#e�v���`�,�Y��^"�M'��P�x���rI]US3���iM�*�z׳�ȩ<��8 p!���E0�h!�f�n�$U��y��*�yk5<�9h  m63u��Q 1w`4'��ES��68!Zw�6b�\��Wƾ4Ү�9���V�FjA՚��L��
��@#	�r�j��~�)!�|rZזaqN��>$�M)��c}UL�����+�\��U��  �!��)�F4��&J���Py�A�P��y[��C�V��{h�oZ�$��%|vI�����B�Rk�n�Kc	��D�e͊:��V��RD:�7�М�REH_����#�b����R�JSت/��`	h�AA�  �-5�� �ó�Q7i*c79w� �p!��v�i�u,8)ts.;  9iΥ���=�@�
5��"���2���?�<
3�j"�TkaA%6Zčh��f)�GB��Y�z��i�<<2�0� "�ITh8�9[ d�ug�����5�����9��ꁲ�-L�IHJ����� ��Ѳ��1UN(ZH�@    �!��4�/!�A  ,�.��J��AX�т�ȫ)�3�te�Z�l91�G��Cg}�D���j?{-e;���BV����D��-b4"���19�<_{�Ԏ��Lơ�b(� ��J��I�]ǳ����7{��9���ѼH���l!U�h 0    !��K@�B5UBft+Cz��
Ϋ�P�_�R�����
N���a�%w��v�a��T#A��uX��[kj�/Uok���L)�v�[n����*9e~�*G�������G�OP�R@ lk��7܃ǿ^�P+�(H��4��T>�ԗFPR�     8!��`FC�"�F���i`U�ڇE[��'�Y�言u/h{ڈ)!�k^��zK<M���7pa�#i�t$W����n7��+�<�
NQ�B�^z���b-@J'��]4!O��[0�2�Ā��5w�Q����Ft��x%-U8�IU{�;�L�a& � �n����Q�(�0h ��I�w   	 �8��}�0��5�CN П<֤�P���uy��?һ^aW�c7+�>N���~GtS��$L�.�Ϋ�i�"`�6CoV���n�5����&���t"0����i��?dv��#��Bu)����-!�{,Q ���i���D5��dC� h��I6��	���"�NT�#ѷ�S~� �'���,!��=u�]DW��V#&-��%;�v׹�?e|(�S[=ir*��ԋK��t!�HPM&*�1���%X>��L4r�߽i��R��I!���4���oZ����y�Ҥm������3�`/�f0a\��$�wQy�Tyk�4��v";w�a�nX�㱐�F	}}L�{��d���Hb���g$�h�n�ŕ#Mw�����*{�Fv�Y����V����v��8Mt�T%��U�h[�|�|���}�\
ҷ�D��|Y_r�*�4�j��t����4�b꣕���Y����0LfK��*0�3��P(b������$� �C�)�Pw}^ͧ�r=-�ݣ�÷��)W��o�Ν���dg�o:��A}�&/�C ���Ό�j�E�R-�Ѐ��`��ѣ�DԤq$���|&u�$ݩ�+��Zz�]�::��$#C?��1��7,7�3{B�=�!sTf�UP��x^�ZFފ���M���*@6�0�&�9�\ȓC�vks�:���L��}lkw���1�R�[2/چ������b9ڇAPD`6�5�"��x���r~�K$)P���u����V��}�B�KF�
Tq�(���)���ܝ���5V�(Y'b{S�2dV��u4����8�`�%�TzC��7�N���쥰p)L}��e� 9�*����O\h�t��-;�5�/�)�y�����&i����;��.��%Z���g"�!3)P��0R5�B_(Gz2�ft\��?K�ކ��s��C&A%qX#"���d��U���U��SX]2J�5�v�{�3�	��>��އ��Y��զ6d|���+���,�4U�D62���D��V9��2,�n�����F�e�ak�	"7�URS�tc�Į��A(�֏5�@b2Ľ���������(��?^�	��)E���5�v]�6<���g`C0����19�!�mu��nK[J�W��b!w�7���n��DWl����1��as���p�����2p�� Ĩ^��s
j���U���9�.946V1E j��{�p.��E�J-8�z`���,8fu2��8���uɔc?�B��>TP@��K`��`NMq{�Y�2��w�<��^���
����A�d�5���GJ�qo�UZBm':��p�+&��A���)����a���k�P5�ע�I�7�������੠;���"��'��	Zի��y��}�������!0qr_H�Q�d�J�)�#>^���{�;��?�{�5C-�:WӾ:֣x�ߓ|�� ,�͔l�-[��u�uΡ[aHKd������LN�"�*Gk���|�`�O;�W5/�R3�>�.7��(8&��r���M[t�A���2bli�����t6��j�H�����*�X���"������ �	P�6�Q,��X�Z��-�K�x7Jm*e#V$f�DJL#�D* ��~�w�TS;�9��]�pL�?�����_mO7�
�:��L�&�I�O��\zvKR� B�.������d�19����aUj���_pz:��*��l�36�k:�P���l�U�L�̨�׃��j�!�\��:�*�05���x�Wz|k�,�5��R��WU���b��N�{�`���Pr�Q-X��2~�`���w���C��_�/n�B�'�,� �G�9�bʑ��5
�^�u���E���������os�sp9}-���T`*��בTR7�ܷ�W�y@�B��Wч�/DZ܅1>���#t"6QY����Y�������3�0��Xp�Na��Y���9P3�i�J�y����O�6k���>O�Hb�o�ޡ��x�wk�Q�����/��D~8�K�!���軶�E��~ٛ�&k�aO�H�f��c�D �L{�����p~��0�FI29�ǖ�7H�qĀ�e=���gE��ځ�UM�&�f0xJGjxʋ�G�T|���\�!U2�}������4t[rp�W֞�x��ߍl��`:���x��e���f�Z�9�A�L�kn��ҐZ�%�Ӥ|̀���/9/'2��H����go|H�Ap��V�������Ԏ�*CY�