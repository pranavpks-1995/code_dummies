��ّL;i���~sT���T�2-<:sV�e��M�-�nji�<L�XXĺ��J�^�d_?���^�&$m� ����TPƺ�{�vzy����ή��c��YiI���u�,86�u�p��x   0yИ����C��G���p��2G�D[��jm�L��8�􋷽�NR�(�!����Ҫ�A*>�l�v슳w��U{�%�aZ���49g�U�D����GR�xcc5��Ic��)ߏ�lz��]qw��ح��M��ga]>�h�c2�0[@��/�	n�`��\ ?DA�M_d�
B<gnD�A��G	;x�G;��cZ�jn=��S�͢��<u�m�������5i�᳢X�!<�C\D!��`�R$��]s������B����l���@�Dt� y�8\Z�s�M:���M�Sk����t��cA�:�%Q���lO��=)zEڐ%��~�YE�+Rj��g���!j�/3�9�8��8��*�Y�s��W���P��c�����!#�k@������GeR~X��9j���������0�䘍N��>�Edb�M&�F�:Y�j�dH�{�� �� -M�9����N)B9�)�_�v[:]����5�D�W3����K��@�ͫʮ�sp�(��3�7<b��R��۩���̰�љıp��0���_g��!L�����b���f��˽7�0W�����D�ͨ��q�V.N�Gk��t��&�&�ϭv*���wbH���um�̉���%⼖}���gx���m�;ݮ���Y-rz2��<�������� ��?���K��Rx���Žl��_J:�q*�n���=|[�.�rz�阆�0��O�X1���I�^N��j�Vf��簪����8g4y���s#$�[�8��˒ԭ�<�fɦ��I+On����h���[���4��V���6�;�ގ�k��s�
[X����R֮gw~�1�⳷����s�%��P�,��<��i�s�����({/o-��-p�~�6I;���N\YeJ��0�g1�Nw�W�p��ELe����<+Ds�?�F�X��P;�� �f�C�5��r�rAd�����\��(P������u�vG. �xM��t�S��8T���3��j�z/Rc)��E��CN�_��7J�@\�7��Gc���I����xtm����A����6c$�y"M��/(����b�?�<��@2J�4��*�?`�����>�:-y
d4.�f׎��Pk�-�0|Hb�T?Ht���A��¹~(�=xK]dG��������t&JS�l��]|gE�K��?��VVS�ۮ��+ך���j:V*^�n�T�H�:f��w��J�e]-��Q��|\��ń9t3�iPٷ16t�ӫk������BgZ�����N��P̲���\f���G���x�P��@��?T�! ���+�L۷��h��@h}�\?(�y�z���P��]v�C_F���} ��LP������W�G�2�˙����'b6mu���y�Ӱ�'`&��s�~�D�4���������`��Ž���@N�T��<����[KQ������7Y��$����/Γ�p����Q�����ޅ�ؚ�i^�+�)K�+1������,9?���]H4���~u�{�}�4��	Yv��nI&���|@��0�J��K��Dx6T@B���Ȕ�H��}W����G�44�O�3��{�V`*�j�Iq�b��}�#n������}�;@f�J��} М^��k�a��^C���Q�Y��W������d�xLd�uq��!���1�2�k��	�GI���ՙ�6�b�먢^UAp\ٿ����l�N���V�Ĭ=�*���ǲɺ�2+?���e�j�e� >!]��4Ёe7v]iO�� O:[v��x��Ϻ��!3P����K�zc�z6�@�P�	ƹ�%�(� v8[�B��ޟ��������_�����s߄�X�}��-`.��ˮ�2�5Y.Ĳ�e�D�VQ,�����wY�+O�}�S���3U�-l�qL����sl��N)ֽ(4�hչT�"�q����sC�c��z� ��q���W�F����fb�4
�S
�D"6�"�h%A���^��^%f�6�`;����*���\���)��̞_�E�L��f&=����>��?��0�2t��Bk�T��]��Ik��}�y%�^-s�l��R�������?'�<�1��޻u���!W�:�g��@��H��l�y�M�:"������^�$�<�x%4����N��G,��!9���x�]Q���w�A��E?�";��u������BX0r�#��b���P�e�焥A���c��gc����͟�T�j�J���|	�,�2�y���s�RG�K/p��JS��6�|�M�`PZL��ܮ΂�j�x�4���D~�)�i��ߦ)�)%�oC�6�'�� ��W�k��l�ARx�lΈ�mP�*�@��� ���syW�n���~7v���M>c�kA��N.�P��S�T���i³�@䔨}[�j�*�%b��,-��@��w%1&L�KFE�̸�ഭ%�b��}����`/#�Cn�*\� ���3�Fua�_cП<�힐���4�.��	PC�H=����qo4=���I\�?@�q����`d|4�#�ЛaA�#0��6[���bۗy��`O$�y�30X@V�n2L�v���IpMF��,̜*�6�Ì�+(4���A?�L��Z����
�����b�.��8�nc�׾m��T�&7�߃������77Q��f����������