��pc�#�F7�z�<rT�Ĵ�M�(����mx%�O+H�u:�k��gn�/�$ۈt�,	j�g��rͰ����i�&O��x�c��a�)X�,�	��F����EͶ�T���9��6B*��D�S1/K-����SݯZ��qf�v�_��3h�"]�9#�NU�7��T�!-��(����)�ct��4Q�J:,}晁�@D�K��'��
��c,��*I��f�t��>�DkSz�꿟�6�.§�z؜��`��8O�H-Ȥ����o3�,����a���@+�yl���ȯ-i��ΡQr[��~��� �����U�3���`l�i�b���[/�h���0G�Q
�n�`������Գ����K�Q�v����$b*<B�m�Ӥh��!A�w��}xR�EL�}�I¨���j�G�N�j�sOQ����勒C����+�\��^����So��
�D�F�����u���i~o%�<����UĦ��Ia���M�[�h�k.l���<����jZ J �q���@��6٩e���ou��[�k͹3��N��78�rC_��j��>�vb�m*@\�]WS�"$�U�p��(¯l�=�_aO4�F�WL��G�R�݄��b�?�`��6 &Pb&w6��ժ��r���`�CZ��`5\ot�R���nS�4XS WL�B�F��6,0�R��y�M�Y�}�w�R$�E��ӂ�Ss^�f鯛�m�7O�Z���,�*�O�wM=r����=b�K�G�Dk�Q�c��h���'opdR���X5Q�st�#�*���
z�S�Y#�L �ܖ�G?�p6��G��������]�yO�p��:���������H��P)�q%����c6c�	��LA͋o0M����K�L��'>���ZAy����!F��� �������hC��z�GX��r�h$��%9�f��8�}�&.i���l��>�YL�~���E�����ʢ{-�a��6�m��H�	I×�i�x�D��lHO&�"jҌ鼼�a��������X�ۛ�mc��s�#`��cz��(q��6��_�D@���sCUZ�:n�m@�7i���q���H�hRO�Q-}��	mi��N�ձې�<�S���< ́A���Θ��pu��"-�D�����,?������0]�XU�-)��\a���C����|Y�n�G��<)�܎�ͪwÆ!eq�<�%i�,�X�x�%[�v*Rȯ�ry1�hR�o��wU�v��f4gk��{z�к����tY��Z��zU�]2l���	9��?�:y �2O��Is̵�a���`|���3��&`�<\�h*֘ohuE����~���r��:7+? �&�=��\�v6g�*������
�//�u��K!6�q  ��+����f�iu\�55�Q�Ԝ�d|�ֵ�1�T*j���x4���j/
F��"Ύ��V��?��l�K�y��ɫ}�"-� �� b�sbI#S@�G��s�~ӏ(����]�J����4�����Y�<!6�=�����?krǵ��2Ny4Z���_D�{�7/���2���]����8<*�zE]I{5!M��q%�� �\�B���ߪ����G ݹX1'ު �)���������S�Xr���h��P��zO����hy��h��t6���d�g��3�&��8���|�'�͒��δWFUL�E ��Z�z�ĩc��ة�Rj����K��52ˇ��3����B�u���-)��W�_R���.8m�W_��ʽ�i�:Y+o�XFe����O�(��.G�V���s�I�!�u齳�<�,�!���5O�5<tq[�)��s��T�
*��*�5'x�
�<2�5u���7�÷yU��0�{�P0���!4$�fcEq���P�њZ�����ǃM�08������D2��y���]M�X�9����K��z��pG	�o֠Zɼ�W��X{@�vT\~3+�j�<ߖ�\b� t(SR��OX�2}�#�Ӯ��)2y��W��<^1��
̛����y�R!�k���ר����c�.3�Q��y����!)Zű}k�q��db���C�I���G��-I�Iml���.l9���e� �������X�g|���ġ�ͫ�̿��H��;Yd׸�� Jc�φ��ɽ6A���$��>�j> ��z�҃)��FX� �&���_����׉��tI��$��BvF��*�LB���S��(B��(�a��)tO'��9�Q�R6���y���$��哅��(�P\�I@���y���O�3��q���en�9D!���|0��}[W��O3�����`yS�W�e�9X��T�ֵ�
K4�f�ILh�.��[��<Uee��MeC|j����u�Eq,�qiVԏ_ʁ5�x* ��3L����E��l��H�+	��r�rT�������v��2����G���E,*�J�VR<�Ǌ�Z_�l�\����k�6DRb�������b��6�l�z�T�N��?���Z��F�w��z���eu~��<�6�1�}�wD�vN@:���sn�]L!؂�\���R����!��>�����l��#�=���3=̬�'.Mߪg�`��!t�͡�W����~K���R`/f-���� }�J���@8Y7>�q�v�(�f2�
�n�J�O���%����I�[�m�P㰼x���r�XŘ��I��T�M���>�K��}��|>��<��:U�3�t1�l����ᮇL���n	�k�!B��=�Qy��M��G6*�+c/"�p-ҡ9��N2\lc?�C�W����A�%�,\���&N�^l7Z�T���h`=�F��h��nN~
���#���{�˱Iȋ����\ֻ^:o�^$~��i������"u!��Bbk�-�FJ��z�8 O����dhgsi��p*2��J�W��h����M� ��s�H�BL\+UGS	�dѦ^��הS��`7�׮����������=�՛E.��n9}�NNjj��\< �xp��l�y�9&���m����xCa���1�x�P�ҁ6�����{r�u6�/�����$��(q'z�[p>�۴���PZL�E�C����i�IП����bī�b��	�+��5(�$�ݯWF�k{�B����k	���8���ގ'G�Ԫ͡�,���[�Gj��R-.��s����	kO�Ŋ���ͪ����gr�5���͸ҹJ]�͔�o��t!B4+9��LB�fc��ϐ���3�R �� ��_ɫ�6^Sd"K(`��O;RJC���v&�?k�n���)rbzDI�[Q����(7�k;�
�ܽ/)��_Ћ(q����|?��zuO��r��e�C[�J�T�"��������h��p�� u*��_��c�*���A�wc���}j�&�r�ݠy!���<S'�v�~��]�S�NX�Qφ^�ʝΙnOLLZJb����kq�n��Nr�e��bW`�7��6�"�Yw*^�z8 �����'�S�'��q�2y�U��J�oc���9Z3A�����=�̣v
�	a�!�<d=�zY's�c��Зn�D�A�����1a�l�#�j�q/�Z�]�%7 ����߶��n�Y2�l++���ˠ0jf���˯�!�hL~�=˝
��4�oG�ⶄ�GKR�ʌ#xmM%�+��P��x҄��	:-{��Ň���y��K��%���N\�|�)E�vd]HSИ��C��� ���SD��	�R$Gh�Sb�(�.��»�X��������B�4F������iSs:��)�G�1��r��ۣ������4�XE�k_l骫�P���U������('����,��;��x����G�P�G��!X�)������'�3��'K�f�0k؟Z�M\�������P7!�u��`��k���a=:	*�α�����m�LKCy�����3����$r\*Sd�Uj������Ju����L��+0���_bi���V`]JlxS4��J����hv+��E6���d����H��5W�Xh��в^;��̴s�E�R���J��]yߍD�0u݈����!�vռ���r�a�$;�8��u�3�^�O[+_8�g3�M5Cԟ$	��vQ��'Z��|�Ʈ~�Կ�k�D:n���O�5�$�q@�NyJ.���`u��GѸ�~�nj)����=�o�*�Y���~�����V\>!�L������D.�r4}ݷYC��]Y�]\�߫�? ��+�X7�F��;-S�Y%�vr*ʐ��,��R�[}n�GCF���=f�`��X1Q��يV���6��Q࡬#�PM"~�c�uG��#4@R�ъD��Ȳ[���c�� ̩�_�5(��ϒ�mr'�k�l�+�sj�"LHz��*w�m���V�`��+�B2t4����h��?E
�	)UY�C�"W�g;T�Um����9����w�2���)����}���uzA�b=z����v.��Z����]����y�s­���(T�=Α,�[�.�S�����j'����6���-�U��Վ
��>͟�6V�@[��ҏ��*Ь���b�A�
�gY;n���My��	��j�>���6�H%F贄��"u��\�1���g�g��2�;��5z,kX"��hg�)b��Doٿ�cW��3[*��Xo�1&ovI8f7�L-��娖��S������旐��o0��6K	�Ǣ8*i��7V٣3����1=����|Ms�Nd��$��!�I�i�����ӈ��E�������*��}�!o�u�� 5�Qg$������*a���~��ބݺq/��M��h�^][^oe����Ff�Z�&�CR�<h��Ɍn؛�o>���㑥�4�r����vnqޏ���Aw��Z��K����1I֭.��bA������2E�Q�E�3�����K�sÂ��PF�r���1S��V"+������\uE+p��)y�����R��o�]�@�jU�d A����|fb[�	�]���QX5���4<!vM��;aR��-Qt�Isf.0���٥~e����Z����_� ïc�E�)��M ~�X���ڱ������HKY-0�/_���_�������R��}H_��'�R;����i)��:�y���wZ�%�!#�ޜ�{)��G�F�Y���: