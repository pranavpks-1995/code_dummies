�UD"ZB�e��ީ&��A�}�dqa��U��o������������8�}e8P_L)������КN���_�6�{��sGV���E��%k����G{5����8�֡�8:��1�̓�y�~ɝ}�L
����$������<��g�y �	o����v���{E������c��ؙ޿A�ٺ3�Y�����ϒPn�E�z"@�wY��oM����	G�d��׊T��,�ϧ��#��UY[�l!�~jGQ���!%�WO5CKGNWDBBC-Qg,.ȍ��7Y�Q b� `�[���,hNU�a&{�����.O�#1d���_7�����׀���g�`��,F_��T�'��1�q�U��C60��>�}�I���="�g�t
����0k��7�h�Ĥ��� >�_^�a0������ڬ�A�`��X8!�������6���(5��_=�K��	R/#�<w��)���b{_��H,�ڊ[\}?��~ҿ� �7("|��-�Ew���.Y6? ����_S�9 Hˉޠ'dIfw+�K�f�7Lx���bn�
`���N7G�'pj�\�Z*�� �n,e�,!k�!�g]�be���NP6&6�>�=1��<E;��L��y`C	q�K��l�y����!<���̇Ux�_� �����e|VB�Ҏ]��1��hJ��]�o'�LmwS���� ����vo�4�ÑQ� y᫐�|��Be��2]D�hGɁu]�(�c��e��