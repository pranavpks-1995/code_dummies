"'%�5�Ț��IԦ�L���L��O�^	t�J�ݿ� �N�g���S<}�R@R�?����+�Ȉ���@@:]�|��֬H�iťc��g��.�v.^3w4��Z5 C={�e�u�oPZ�� �_~؎���XA����H`�����#�'	R<;�pvR"�9˔e��,���wax�X��Cwm�K
Vڬ�˂���E���|i�ũ10Z:,��v��1�;>���I���'A���n)I5W���4v����D�IG�^jT,!8=�3��9�6���|�
��ts�A�G���%�}�=7\���)��&4����8�X���q���r.�T�gs7�D�xV���j"�C���,�pT�$���U%��������༫�) ��2��T��J��V@�Xy׌�'�l��⁂�e�����./�(�H&=����@�   � �f��H�х��B8��R��f�C��	���N�q�l��x��๪�%璗b_�5wC�^�3Q�]f9�-&(�7�����gi)�]���	}W]��pvRђ$��:���%ʊʉ�#��H�V�d&�L?t��*��<��n̓l~ez���ll������-�����{��Ɲ�e�m��x�� ����!�бU���~��:��_�د�*.��L��C�u ���9� Q�  �  Q�*�8]"q� �^޵�ۙ�!���i��<N���S	�y>+e�k���p�A��8����Di"������!d���!˖zG�M:�*	9����>��D8|؎�t,���<0�KقW�ШZT�9~�-oJ�!6&Ñ�X(PP].����%��yDR�$�}��c�d4 C�Q�Th|͛�G(�Mj_�t�툰���X�����"t���Y�Z���s�
���;��9�"��շ��XRW�������5�)�)ez�a��:��`6ޣ\i��U�q;]�1��Ì���
��?�;Ōq�6�X�K�q����[��*���nb���<S��y\g��^x�g|������Q�Q�/f7�b�W"�s���QĮV	A{A��q�9V�g�c6 ����Zlb�=��T4��]�8��_P�k�-����XuEU�HD�(�5��S��|��_���q2*����T2q�ZtE��A�G엫�V���]L�ȫ�=z�J#w���/7�������K�ڟ���8^X�����r�GOGb=:{?6�7�y6����x��X��U0uU���n�A��; Z�P�t���=�l1c��l��j�x�[8i2!#[c��oDgX4)s��KUȏ�����=�A7�L(���l�Eܿ���� ik�d��IY�����]�Ρ�;Ǖ6����i6�����v]sz'���� l
Z��⪖�؊�K�t��(&�L��f�96���R�^��R�bD��_�O��!;���\��'��*Ax�ܠE\++���ږk�\����~!s�^������zU$�:�
��-��>��V!��}TƏܖ:�P�2@�� �h�Iq�8���#E�9G�7�2P�PFƳ�hc��>V������Ez�թxc��%�8�(;xL��D�^Z����x<YeB�?E���g���1��R���J�B?��=@�d.>E�Bg���H����Nߖzx��D�z�FL!*S�*��D�:�����6�wG~(���u7���,kNC��/Ex�����&c�E����aKJ/6������Y~F �K�-�+|�\�	[�8rJ�R4'��Lk;5h����@*����S��e�D�~<Th�4��y�@-���^����}��؍��0�\�~H��1���,���S��uTއ�`3$-LAܾ���	.�	%�� m��}��m�_�>lp�`��@&C�d�a�[ޙ����du�P
�sR�J�f}0�#3Ƌ�ﾺ�RGOO`�G~�F��,dv������xѹw��a��}ɋ��