,杭�bS��G���+��|�'v�}��EW��}�a�!�ԩ��D��D�о�1�3d�k�d��,��������K�y젥�JO�KN�vJ?УAׁ�   � �B-W����Ã��� ��Q6�GV�	H܅*��iJh�F7lx#2��)��ǎ4��/��\^V�w�M�T���S����h��0�W�7!�~���C �<�8\%r�Gҹ�A�mk�+�+��늴aQ����'�r�������ďTP�V ��ؕ~��ֈ������rA��i������K�Y��u#��)��]L�כ9] �����d�=7}	�`o��Ȋ���hh�NA�������c��r�� H�47#�ɬɆ��_0}$� �As��ۀ	��!C��� ?�!���V�����;��@�d��%n|�R<�.���!��D�rv@�>A΅_A:����L��DN�*ܲ�'��O�2H�a��Lz$"v���S�����C�� �t�#7#9It�~Yu&<'�k��̆�ۻZ�mS��R�@�$Q��P�9��F��x�^Pha�ƓMf	��E �	W��������!���҆ ��D��-D��W�]y�ӻ�t����*XO��uY�1b_���Q&L�ԍ$���q�

i���$?�,�:h�:��������e(����*�3(m �b�!Q=����m�t���7&4y˵@` р8!�Ԟ؈�Ġ�{������y������0Ìn@c�S�ދ�VJi��]�_�ưH��N��v�[��vb���3V]8�������pn��p�=?�b�����T��3�}��T[�����n�&a� �V�ۤ+)Yh^�e@l��!�� iA��*e�p�.P����q�i���b&7L�>^\l=ϓfT[����:\�d2���"%���@B����6�R9����K�g�����:�!��5������^u��w�Q,���M$�T�A�Ȼ I�����no/�`i� �!��Bb Ȩ b�	D �F��v��Wy�d 	�R�n[�YK��J�Q&uT��Ŝ%9ȩ�ro>B�j�w����,��x��;���?�'dR�INt�xP
���������[L���iRC>�i�~9�y�	�|�w7i
�\#2|��hk@ p!��5�B0L�l�Z��7���Z�� �����4w'\,jhIP��8�uw��蘮�=���\�Mڦ���%���<��?Jep ����]�A�J4�8�7��Gv��� �CVY%��c󎻂��tuz�$m��RR �A���m�T͚99�"   �!��a�X�H�"
+�*�e�h���1�m�!R5ү(��o�9T4~9�:^��%�\.�>��H ,��u���H�Su`�Q�z�a�gid�g�G ��%��J�W�E%��?Z�� $�s�>$����h^I!tUR�
��V�.罭W�x�d��,@ p!��)��������bx-���Y)�p����8��\�W���j�Ur�RN��h��w$!) ��bT��u�\[����G�Q�1��Տ��~#&`gy��*u�D� �@('��V�����o�,a5UM��?zњB�#0.hy�  �!��MB��B���Y .�ŀ�^#rK���IN��!� ᩛ Y��U��4XL��x�8f�H3y�_Fq�-���+���턩Q���&p][�*��^1H�xѲP�ڼ9�����sE��|��&J�
Kժ��k&J��T#�'�Z�	u`V�  ���� �+���  ߠ��@�� !K
��P  �N�	�   ����W�C���VO���#�.b,��8���H��v���黯�����c&�����;$����ؾE���o�N���?�c�v���[ӿ���~��Q���i?�8��2Q�F�WҪgh,V�#::��:�B�DP��|�f"�n0qT�	�!P-J(m�ʁ(0͞���=�P?i��M6�ё�L֥O��R/��L�x�Z�3�~��g��ܾ�dn�p+�&��Jy��B������Kt�o����@��a"/Ơ�`�t���K�6"F���1[�+g\os�η[�����T���}�c�X�>B�t_���<�I�x�;�aN��>+gR'�p�f�\m��-E+Z�t�|!S���f���~�>R���t]�`�2������h=�����cG� ��+F���(�u�����o�����_�P>-$����Rv(l+8=XTkH\�|ތf:ea�oy�?n(�SBX�Qr)��6�Y��H°26����9����� �5��G�TE�#b�su0�	]�oe�٨M�QV<E�@� �#٬[i�3@5}���MNUh���Q�E���C�U\�T��"7��w��^��I������4���v�pJ��p�z?��A�)��G�cy���vRS�W����, ��F{�Z����֟�	�_�٪�4�o�}�D5�a�tDL$i'��B�T���fB��6�R�[�/̲4/B��-���dW?<p/���@m	� �+�b�q��
�3ךA���WUt�������Dӧދȋ-]1�􃁠����ޛ�#�U&��W��7�1��8I��s������mݽQ��� jB-^8c8X(�l���B���n����A�p�g݊��Vx��l`_3�*7�)Ȅ��E��h�a��M�T�{'H�կg*S�Gא�wѱ�\��s�z������y"�&�kZp%��Mx�+�Ƶ�z��3���+�eD�	k�~G����Bm�N� \���浞����ٽE0����]�mz�m�{v��r���j�*���Г�$������ѷ�P
θ��#�;����Y��HtQ�wv+P��gm
����B&&\7���a��
�ZA�D��+e;@��xe�5�w���4f6�z}�ođ;�/�y�HY���-R�i��!�ފ��#g�R�����D3���ϗ�D�X�c��1^�w���,���O�@��n�U����������ir��ߎ����)��+��"�*\�(�{����;�C��9�"���2��Rc=�w��O�ȧFD*e<1��z����=-bu��P������4m�����8�IW�a�"L�"�%�f_�ev�̗൅��dO�7^9����CJ��a�=\���#f��HX͵�9������
�D�b��d�Xw�r ���i�d�����w��MU���i�"2��M�g���LJ��I�h�i�ȴx�xk#-�9m��ҝ�evpK�-=ͥu���Gؔ��m;��*ނ8��5l�{~(��S�YU�������T}y!����s�(נX2#�^�YR�ڒ]	ԭ����@_ 8����"�$��Â�?�kL؏�IgV��|�0��;*b%����%�Q��u�}��Z|�͝�Q5b0e,��i�j����]���i��;�.�A�f���)��3����@���k�<�a���y��a3w��l���*�[}-ƿ�?s�Q.מ�r*�۱H��B�����>�}媾�:����hC�UC[F�ܙ/�'IѾ�$������=r!��5�����5�������1!�(��E4D	0�q�Z��s��Ln��o���k4�}�;
tHE�[,����?�0�%�^����Q��F�f^>�i��@xM���;m��kͼ� �2�␞���ib��Q4ٍ�=k�w�z�>�uZ`�P#���S�F�?3�E�=�e�a�������Ϧ
��lx\��z�?�:���9�z[�_��@��EV�x���)�1ۥo�+���W(x:m`@�`�wՋfx ��G����Z5+x�Z<;#�
� ��-B���py?��!����Di�\�[���g��lHo���)�&R=���r��,��ď;�R��ӣ2	gq��;'��N�{��
�o�����U�B����h���ٮ��F�iPL������淁���٢a;=BV���q?�A��g�Q"�R���!w�122%K�� ����i�V9[b�4}S�����`LA ��I�F��J��<�s�o��V�k��v�-�D� b��>樓���\9�Q,��-`�c�X4��Y� ��ƶ�� �B�,y� :���ٵ��$z6�4��2�`6r�x��P��S`~�ȋ��kWW�~����&k�eĦ~�n�پ�Oڌ������Bpvu-x?�?`�ہ�m���=�Ȼ!����GmJ(#�vض��qT�`?K�`�3����ȫ����zy���1A�9	;�2�:����.��g>�)�^��<����6��^�>[	d�x.���$L�Bh�c�R��������֎����S��{X�w�],=�z4��ڌ��Ԏ�陁��F��Z1�O��#zl��B�xx�)��Ni�XT��.`��r $��B���/S1^Z@Qr���}>��]K-6��hbӳ��H�t�u��M�z���w��0F�}��ʻӤ)�%@�i�yΡ@}���x.��8K�3h+"��H!��h إ��n 8弧�W��H���3��=WmS5g|�bZN�ShX9Z��FҀ