����m����J�'e8��� ��|XX ��o>݄�l�B�Z��V�f鮣B�\H���/��T,av�F��YpQ���_���Yօ8BP�ϛ��kp� V���#�|��w9�7�8	����������~�|%ͫɘYGH�<��ݳb�Y�N^����.����U(�A�CBI>vNMFL%lG;���0�'U�Ae�8A�He��tj�yȆ!�i�u�R��!"�20Q�i�?���]0��79WIݐT�?�vsU�|�=�G��Z�N��w�S��q��e0�X�wYwi�4�^?6�g!�h2-(E��81*kQŋ�Zex%L?��zp���>�ٞV��W�6h��N����J��!�4���֯�1�=���.�6�����p��}�r��~y�s�zQ�r4ͫ\��p��X�R߉�)_���πg���~Jk�z�X����ds��X�i�P����D$�"í4>�re���7`��Qp��b���	������5���X^r��aP�mA
�/��Å��O.�Zm�k�u��4��A��������-)R��V{j��29�����U�1�*5�fd�6۩Y�*Ap�j4(�=�ݺ�|z�2� 	��(B�@D^+iQ&�r�7�2c�c��C�ɹ]U=-3�VK��|w��6�L��~��,eN�f��![g�����Ʋ�~FYbiZC��ʡ����c�H�q�.hIB���v H��<se}#ĖN �>��V*W��B9�j�M��m�E�ɸ ��`�5�q{�샰	M�-[�����.�Z"Ж�"�5=�#n�Md�@���Ο^֩i���2-�.���t�B��d�r����I<����0��ŧ1l��*d���������hh�V9��O����݅!u��Io�&��'�g����� B����JƄz�Fc�ٷ��3h��k�ߤ�7���p��9O3Y!�V���Bw��!��c?�_��7^�=kX/�c�3��U�êW]��k26��Ìѷ�\���n�3_�7n��oT�oͪ�����Ys�(?�3����6�ה���h��.�a�ǎ;��x&���Zv��qZߊa`��9�8:;�}|.�[UW��<�!�?.yc�֯k��0��1�twZ"�v�6���K��!�L���*�<߱�=��2��"g�`�G�ӧ�4��۫o���]��Ͼ��eHi"�檕c:�dLp��-+��$Ȧ�<�c���e����zOB~y�`H�X?j�3��H�~�����QY�
�����<�<�-D\Z�pVvY�t��[�^U�W�\-����?�0GrԳ�J|�D̄�/	�>b�1� �Al��`���3���m��� m� ������LBs���b�y�J3�������(�B=�x$
!��2a�yBA�cp6��s4�w�r����R����H��č|sY`�_�rMς�δ��5rF[��1dh�b"�9?<�,�;�N��z��#��	��F��u*����U�~m
�6�@�G��2�&s�uﰎ$3O���p�ǚ
������%~�$L�0u�����Y'����nZ�<�>�d���9�^)�;��dh]����Y�R���yԘ�����Q�p�x���>�DE�(-��� ⋮��<TF2��8��\�f5�e�B�o�Ci6��P�I�7��v��6�N�.v�"�c�T>��=�W@"�αdS�\x�B�$&�:ow/ȩ�@ٽ���ʌ�X�^�P���Rk�@�".�g
<�'ȟ��eo-P*j/���o�6�Y�Cy��g�QCă�Q�`��J�y�� I�9`>��Bd�}g�p����\#9œ���_\<�ޕᅎ�k�Rً���sԻn-���ml�#��&@)�!D�=���*��6�B�D�֞C�WH��l<��\F��kd�|p~i�(�#��D����`.A�A��z�!����=ů/��B�WzzP�ٛ�wU2���Vx��{����i��r󬨍4�� �R��β��lk@�H3]��bhM:ur��%��{w?��{�Ē5�S�	z�7��рjJ�_����L}��a���ȓ�<'�U�����C'��=�8����Feg�o��hu�p��'�k�Q�Z���̧�'e9?K�9�0���8�)��:ߏϓ�V:.So�7O}�U�(��4D���u �CJ��J�P|�R����T�84s����4�-#u�^c�����..I�J˛��-eQ��=o