(Q�Jx5nb<Nh}���A�а@��e�"�O
e��\�;�6"���?1�������tO�ᔐ��Rl�Җ(��n��}��Zw��^Ha��m��.T��^��S,�$�i��(�I�I�.E�F�"%z,�8��Y�-F]�Ɍ���]F��V�;N�Ҟa�I��@�݂I��yAH�\��Q�{5����s��|G�Ұt���N|�zb�rp�k��H��V�A��q�>��<�v�����sщ�Y���r<�o���6�e���K0R0���o'n�R)�4����r�Ю��>�"�H�?l�m�I(qt*��:�"$�}�z���U�Һ|#�Ӳ�X�<�2�!�s9���w2�r�r��2EoB�lz����jM1]�!��/����`����)������p;D�*0��U)�XNG��7X�y���QMY�D,8=&��o�\0o��+e���6�@�@r.�3�tʲ\U��r_#��+M�<���*��B��d�{a��{��d��ضƌP��8E�Fi�H���l',��|M�7e���O�
�%'��@�������3���f��8�̷�*�U`a��]�8�v3J��� !��i�~�M�ߖ:=�۸1,���%9��,.���	�+��*�#y��`�4�s���Ȭe�rU�V$!^(k���sE &L^����K�ʢ�#�Mf�6���0uu��8�P^a��k]�����ȨD�S�p��m�9)ȥfA���_d�i��t)��YRJ���泰�lj��_� :8�	�#�rD�_���*w����>Goҷ�"�S_�5���n\����0W�i�X���dq�0ʺ� "qݠ��\V���*i�Q�������]�c��1
�o���5����Àz>�w~����N.'C��RU10VqG��}�j�t�HO.C���G�N���1_|/l�?lk]��9]��%��0o�F*I���u�F��Fw�v
��)ݖ��;��+�5�/iv�*�}��
�_����e2^���d����oѰ��?I��QǞ(ڡZ�+�	�w]��쒺9b�D?��  7��'RW�c��+�=V�:���٢ȅؚi8H*�jA6�{4�=�Z^�k�"���\���A[�?�i�ҕT2:�}�l���?���%��W�2�Ey�{֝���
`��kk�s�����gt3^Y4q�T����F�iQ3��z��8������=��%�~��3�$�C�R�x�4���~���.���(J]�ߥD{�niQ�>������v�m������I������b	�I0��4�����+;�^&�@n6Z�B5�����Vɻě]����۩�Y�B�?+���R�CB/2�Z�`�DN���<�j���V�S��%����#�Hyw
��ⶀ~T��u�4`5P�˭�f[��T
��U�� ��)�H�)�"��֐H=���ȉw�Hq�:��
�e�\4��#|jr�NN�潙<�w����#��{
yV6����2��Ƚ;�O�f�qV��T$V=�B��K�b�v�e>�����p��yc���R&&�A�㳹 �z5W��L��+�G�w'��Ә�Y���'�q�m}�����;;�bL����.��C�����q�"9�B�>n�����x���B���t��Zi�;�g���F_�����l�RQ���b�Ck�x�����勎W����Hն�I�l@l��D�C���wF�VP��t=l
;'���7�6�<��D�O-I	+��\WS�Jh{����ѵBsC�a,!+��膣�ḡ�U~7�R1���i��nqgPR;�!Q�u#ܯ�t�󂤤1�8����tJ�������]�f=Х:�>'��>#�P�s+��ȻJ ��z����!S�����_��.�t>�f�t��X�	^z�`�zS�o�*X:;@�����aI���(�y��4���j�戬`@�����)qa!����9�*ߓBV�&4��xI^e��i/v׫�誖�M���o�w�	��6-�������ê%������|@y���wSIH����
e6'G ��%"��ҟ�󚻃�dӜЀu*%���W��:�~Z`����LD�D� ���u��Bt�H  l ���U�r욥jĦ�@�����D��nO�����.�հF�X:Fq��6Ph^x��i_���(#q�j97\2��"!��o�
�e�8�nȗ=&0.�˷��a�}8�.��C��Ʒ5z0B�R#��	�F��G��3կ1S�Q�J}����qS�"��T-��C+[��tx�H:Q򻋋{j7��
C���H�4Y�d%3���@ ]���5�7�R�67���a�2��{.O&���-x�U�?Q���U	���M~��TP��Gn�qe��g�7��G��LV�b�-�̻����:x��4�U:����5Y�)���^r�^��ZS���2h���Cz��:��q3
�f�s����b���a�XuE�楘�N&�?E��?�X�(�;�K���\9R�ʹ5K�Q*~N=Ӯ��ʲ��P)�NY�>e��T7p�G�>h�4�X�y�u>&F��9���U���Cl/UA�zI�:�|�"4o�:�7��/���c.\bzݯ�­���F3�]^bt���_ݭq��o��Ao�Ř�`Զ����ɫSG�NJ�JTm��8�h���X���.�����(�y��vxc��5��+P�<%/���` !��Mp`�B́r   � ���u�sر��tև�@����co�E�o ����%����F�c��:���|o9{��^��%�p;e1z�A��P
�:m	)B���@ڀ����"{V�f)�!�AM7��n�l��<vb�<y��^��)VL�]d����!�ȸZ�p���5$@�q�W��$�}�٢	$��|��ܣw��T��8z��y��ghґ[-�1s��������� Y�؝�{n��zPц��R��ø7מ������M��	� ���"���:1q���6��)6�p0�)�����|���8�a�:�� �t�����{�Nq[�C�ӈ�����^��� ￳O�AA�$�p�]�Č�*�24C;V��r�S��ޚ&p7���h�/�zU�§�,	b{�bIVEH ��ծ�.�|��!P�d�^�-�'����isn���������`��������y.9N�Ǯ�fԟ5�7,�\%ӡ�� Η+������n�;��+bE�VKٙS��˒/���G�����> ����:��.���&M&DP��́XԡYU��!�E��x:̿��:O�T�U��:��}��d�V��l�Y�N�`��tuiD����/��W��~�\�$(�Ǽlݙ�!�x0g_�N����3�kC�d�����;wC��Zo	n]!!L#����Vcgp�c%��H�!�܀<��/��Z���AW��   O ��-����"����-:���>Ӗ�y!t��)�t?i�C
b1F����=Q���ϝw�(�!�Q1�Q�4��p�G	�'@{�bg<��{���*�bw�S��;��iل�й,E1��.;��9:�PL.�$-0�ٺ�R��ƚ��2�*��ٰ]����[���$@���/x��$�@�#F�*z����Z�IG����D/�Ֆ�Cf�ܔx	�3�SA���-��ӟ��A*�Ҧ��ѕ�=vs2���T���+o��qY����guB�B{e�Þ�������Tغ߰a,�ZE���>�P�����2��6�9��ȓyV�^ӠЁ�t�yW��I���   	��(����C���e�[����1�`��� �S'%,�~5��C`�Z�%q�@T�,Q��Y`v�O>�X<(X]G��v�-�����B�7x�}�j4�z�o(�gz�9�k>���QŶ�#�m?¬(�wΘ�)O�P��w��C��a�>����AS�o��,@������Mu� �^�h�|kSݷ�D%����n@�.�"F��]����U��5W��
�(oV�iU?� *Q�#��㵟]��XH�%���E�,_U�U[�C�h��
n$;��T�_Y����g���.܁7A�z�hIP������E�4I���؄6<��Qc��5��c�������i��3x3��D�W�G�앬�t���;Fu��� 튏G�e���W��n���s�ŝ��]翙65h����5�B����8���|���rYA���n�a4��������p�h���l� ��[�_�c]�:d��j���n�D6-���Ph��cY��C>��qvW�q�0=��6�<RY��z��>;8����H�ؙ���:��\���!��n?0�hϾ��V-�Չ��ț+�^�`�A�@��jFZ��s��'v���0�+Y�{NX��3Ɩ�5�7���r?���M7(�����3v`�dI���O���X��n:o����ڃ*D�N�F�χ���DZч��G=I�c��dgu?԰\��n�b�Z�s�㡊C�,�=j�	�Ք [cSf��t }��d�\�NA�tĻ ���D�/~���;M�0��T�EnR~x"�͌��Z��)�F��y�:'*x R��P�	��1]�B�JqX;\�@���J���UH��H���1'��c,3騻i�ˀk���T��}h�r�7�?�az��iM���gCWF�~�[,in�"�3ɴ�c��!�� b��4��p}�$�Y��R��Gr#dY(ʡ��P1%S�ob�6�-q� �#�3@�&3�^R Ng��4c[ �w�H���_u?���d?�������\=���c�R��;ND� ~D�D��5 �q�	��1F��<Y`P{�G���()Zj69.�['_*w���a\��5./0�Z��T���ߺ���a�L��,�LT�mnYv�C�n�U��4��� �6���Kt�<x�'�
6�����˖sxh�4��J!7t�K�Q�u��������z�v�8��1��//
ԥRÛ��rs �PK�.et
wW���A:9JVy�e%��}x�Y��S4�9��ь��	!О~.�;5�RF$�&!���CE�Qj<T�)�E�/���R��16�6�M��b{��hZ�|�QB�E�o�G�����G���9'��]��u�wЪ��d�i	�WUwEPY��t�|�m�j����g(mm(�T�����g`�� O`�I�	鶂iH[�D*�Uީ�zc��I�7����v�=
��M@+�#c���2����j��7���t�e����`����>d�d�ouiR*�=�ng&;�~DfV8�q�DAQ�u�
}��:��}��d���϶��{�F�m�Ԙ���-��U���SC�k�`)��7�{UL�K˭3��W᪝��U&כ.�����2�ɷ`�t`��;Nv������F��<�j��� �	K~��K���v�C�P�l���Qv
{)��4�O7��f�Bš�]���8�ܱ��cGeO�g�A4�\'���sS��Wv��{�]�!����#�A��ubM��W�?�²�6���VeB֒��ß+p� ���R'�C�.S�A��?Z�Xo���swJ����o�Ym0jD܋��Ú@ě_��3Q8P׊<�㊉��p���p	���&ߪZq�������:͕��d	%vU�W�$vOJ������=�F9U�������̒���-ɢ����s`�x��@�˥���r���=�/+I�(2�&!7��jot���MZ��}G��.`�^��?Rq���zR}�	i0�;I��=�4�U���$����bU˓ֲ�sŏ�!���r ��"��� �s�gК��AE7f��2<�%z-̏1b~2�|����`�*�#
� ֈ���Վ$o��XF�	�n�+-D��?�]�y�*��e���NO�˄�����������	�5�'�On}:�y���Q� �[�*:�#�h�~ڿ��qh+����CQp����9�}qSg+8KQaJS����@���3t6i�Q{@%`��y����;�B�z|&�ɶ�F)$�mq�	.s�U�DA�y��}4�q3�a�[����^����H|!f�0 �
ޙ����Î�	����性��o3KNش�����=�t�
N�&xm�D��b�r�6xo{
�6�hA���F��q���+����,khr�wm�m����l�I��
=�\�.=*�T��q�{E�FihُN8��!��G��أC�l  �b'R��c��&�@�
�m�;3�Wtp�G�6:��L�M6's�w9Wm�����S��g�@@A�0PKx����vC�7�7�	М�4��u(8T����K�8�@i����PXo}��ݙ���H������S'��M͈�>L*���%3Q�f���%�2�0���t���3r�59P��F�!vx�j��(�mgV�5ۨ�ԯ%!�7�C.�r�
Yd�Zb2���&S;�2v��'�����o���Cw6�����5��3�j�F��L
�,B8	G���]	_&�}G�e��Q�|A�rv�<��U����~�ӹթJj�O���q;w�H���ͥv=���w���)��N���U2Z�U�U�H�E�4`�9C��.֕}���(��z��C��@+N��Yip�(��έ��9���v�����αo���m@>�>�Y�!i�*3�=�b��2����X1�֒������->�2���pB��f恑���&���:��Ce�kRn!8��yt4�o�`�j�2 �ѺT��`�0k`>�?d۝�7��厪d3:kċ��EG귿�l>�$ �C4z���3 T{N��q*��T��QG؄�����Y�l��F�#&��&���x^�θ���^Ẕ������I/�\��U����vm墫F� ��.s��0̼r�j��Q�o�� �w�����f��2�^�!��83eyZ�9J�u��,� u���I�m�|S�
�g��e��B�   �&�U�sƏ)�-�����N ����n�E1e/	H�!'���'��+��,ؐj�sUo	������]މ[0G �o�@k�i)fn��S(KQ�Dj@�V2�K��=*��_珁k��{�\|e8�c�p՚�T��t�R7�nٴa(