��L��"�9V����܌�
��
�I�xd��2��Գ(sB�Ҷ�����f���Y���J�>��⍒H��/W3BoQm�4DpQ_G[!e�P"��R��"�_�j.��k>!�҅�1X��L⬺)�`�h��o�B�שh3A�k�W��2��f�)�2�~{�k����ȅ���������X2���)j4>�N���WĠ*�m�@�b�a�Yc:p��`�uŀ+gզ;��n �(������~3�vԈ�?�����%["��g5��I{����ZNR͸��X៉����Gs��m�7dxz��M���`��I)zVe2�u�c�l}��<�+;xk�k5�`K��C���pR�#*���Q���}�B /�g��q�<m5�<�WO=GW�5|�Ҍ�xAC꥓�v���Gc�+k><pHE����Dsd��{���4������YN�ت�	N�@1�%������{ET� ��~����+�Q�鐳_r�yV�rn��G��!E�NIP���D�L���3�gI�]i�_�}yD;|u���RmQz��!�V_���O9�w���#T
�^}��oG�������2�rm]b��&��Il$���4	�ȓ�	G������8!77��

Ҝ
m?�l����"�_`JM��C��vR�dP�G��B�Ürɱ��gW��A���L
6���^��IV�-�6�7%H	��ٶ�avz���H �}���{��͵�Z���}�k:�$�"���#�>L��R���ї,�w��.�i�6�*�嬋+qG�S�h����=t��.=B��'"6K�A���F�qV����-�?��v��/ci�	̝�R��6ɔ�n�J�5�_~Z�D�q-�[��)��
���̝��,���hIΛ÷�ˍ��$@h\y�Ng���v����5H���]C���s��t�\����U��o��WC�]*[|��Yey�r��CH�6]�P6yo!���G�_��rzѳ�M�$�Z]�C�G���֐�Qm�c��X�]��X#4�q[6P�[|S�,P+��N<��n5�4�
N�¸��������6�w�<�5d��C?����{\���i��(�΢�����f�� QY���]w���-�s��;h��6���F��>��e+f���*�E|���W�h��<�|D�j��xJYab�x�{#	3�� a@�c2ޛ�ȕ��7y�nz��vl�b�*�S�+����(�p�H=�2�G����	/PV]�-��B13������b�ER"Sg�u:�i^��'c�{<���N����yƼ����'#F(~�(UzA`�l�߼�v*�b,ϗ��-���%���`��S]�C��[|���8H�s�+�K�%��Mb� 2?�����B��p�^���k�w��=��۬U��F�}0��}���9%��6J���X�r$u3�_-�%!�Y��MJK��Q3�vtc�tąOmX�EQ�  I ���U� 44P�OS��2^pJ���X������j�s=�7=�^�@Y���m��ӷ���N��YU7A��M(����$	�f[�O��#m5\�z{�4�Qh�b�-c��B�E�+�w!�� /�0�����H��ra�~	�^�9]'g���zF���cv�"�%�E�[�(PMh,?��X��*���s��1l%��:y�e�lE����:�S���b��	N /�Mz��:f���D�y��̾`,A'y��B�0r��vs8�ʉ�1����Uc�P`;1��d9�ze�Ѓ�f�<��ڛwyl���-h�b��Hʸ�]��V�x(�*ox�s�N����J�!�2��� 9s%F	�m��;�O5v�i��ח�:o½��	O����MM�G���s������:�e��z	 " �7�}H�*�bب"� ���7�D��i]�Hk�l�Tr/"�4k���W�)b�Q��+K�8#�`�[c.EȐZ����bhS�k�MԨظ|ى���n>�|�#�7`�s��q��x6U��%�:|���k���-�Mu�����39N�Y���>�:�⇭%N�<!�g�����N\g�A�/�0�̺+�S�Ļ��%K�.�EgW�+Y#� �ٌ�i���
��ɾ,u�[��y�d�(H�KP����_�C����eH2�����ie?Ѽ(�p�^{AL�W�pp�b�-~t�ʄ8��Q��V�����#l�q�~��!���K�^(4I��X�Ǒ̈́�LϞ�Z:Vl=�� ��X4��qi��Q�>L�(Em��߀�N��S���F:��4<��d�F��c\��-S�;l��(�h��_6��>ra�8H�Y�eht�����[e)��R�����'�_3��ۡ���?:^�s%�1<����ɡ��w	V��i!�;�*.~�w>���� �� ����@%�B��#�f�J(�kd.$�Ẍ~0��W�z$�4���nb�=��2>�U���?E�f��%P���Қ25�0�\�E��@���5�o�g��A)�ע��WB�r����Z����\��O��.J�_
j ��T�g�>�˫�P?gĞ�����l����bWB8FѸ�����`9˕Z�������	B[}���4���������2��RoR� y��to�$z��:|����Y񺮂���	��2����%�r������\�[�����x�g^|G�s[�H���X���r�M�������ln�Z�0��n��
��X@�4C�c2�J�a���Mg�h���-턣��G wN�����P�G�>���۟��N���g�H�=���n`�EA�7   9 ���u�$*�ǧ�<!�bM�h��?�<���r�xy���Ras`��?�g�	B���\!�b����=����4��el:	m�#�P�1j�.N$-d5GTɚ�wh�n9���D�s�foB�A������g��FED�C���3�j2��q��p�%E�ɬR��#>��
�B��K��0�3��_�`X���9�q%�� ��]ˡ�o��:'�1��	��
$�@#!?1'����b-͏w
�+������zJj�k���
kD0H_4�t������Ά����h̵�;��.�Ԇ�m��$��Q���!����÷���E���!���� c%���k���W2AQ�zl�f2/á_Ǌ��%���9���vS�fД����ò�I'N6����+sa�j_g��/�����Z�2]��Y���c�o̠���a�����B���ߒ�4�6'��#���R�x��s�fR����Nߝ�)�j�F��Rh�*��V�.�Z�ho-��Lk"��o!�O �Z���Ζ�U�3�_�\d�]��֋����G��"-��%���P���C�G[�[ SU����y��7�����Lb�#��w��4wϝF��E��kA�;�>\WIL�gɝ�m�̿��!��r��U�������M��3b��>��U�ܞZ-<��QK��P_�Q����!I&U��!(�Ʀ`�]�Q�
=���ąw���!�A��+GH������W1LA�D?����qX����O�ʚ�+��K���'Wu�{�,}5���<S4�p�W�s!�`Ӧ��}�{�	�5K�ʬ��5N�1\�{���8�����������z?\�W�m�����j��+eʍ&��c��=��>5Ǚ��~:S+8ɎW�.=J��ɝ�o���Vů��0T����QY ��)[s����R7��7��V��'���Ȋ�*]��3��@edª�(_��_�t1�#����n���X@�A�O��I�p���0J��
�I�A [X���7{��ئX�2��(_,H�AY�.{p3T��Ƃ�1�����V78�5�������@�7@ ���P�_[ �P�:SV��:�j&(`�AoU������U�&�W�C�=wN������Ά���vY7��LB:�N��RL�jJ�O� ��tt���`���R�+$���lD�
����	O�B�&���%1w��r>c3�bI,�5�
b�`@Ud*p8I51��
�����^���R�gA�Dذ~�Z����e���&��]��|�F�7x�=
��{�Q^3�-2~)U �C.��   & �"-����a�D�iPM����7�>�L� >�ԣ^��HA�x�vT�DV�D�Ӆ"u��D��$w���ުY��rH��V�IiN�x@ԖTqr�����x�=b����5�
�|�Q�v�q`��(��)�s-��i���3�ɞ(�-��L^���3D��������͏Xf�wp�&�����e�h�/�