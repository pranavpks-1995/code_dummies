�K�wG	ЊI��B�k�) ��&+a�P�a���@�@Ɓ    � �"-����LyE�Q��8��Gݷ���2]��}�i�[[����p��?_O��S`�nX+O=D* W6SNA��!+�s�#3p��f�y��6S^3 L�4yt��$H�z���>�7�(S�����WFGt�7 �'�g�%�Q��,���w\���� f���@�QiS@�|���ɰ"e�F���IiL𣘣Hv��   n�8����C���dQr���(	�:���O�V��V�)ܼ�U�&������2w��L�B���b�8�e`3�vSx+�����v�	�C.� �ޚ7J!~N�t�s�m5�M��d	[�xOdw(  �d涌o}����J���[c�ZZ�g��/̣<�`q�Lpw~$1ʣ�	<�_l���m���ts�L�S���D� x��O#d��6QkUby ߧ�e�ˤ�\"����tD%�ܞ�)�Ǯ|��Ʌ�Ap�Q=nЌ�x�g�_ڻ�l��P��?, TX��*����^La<�i`��?SDcN�y!����sOx���kE󡩚:�m����`�����ͯ)���^.������+�Ɓ��~r��%����q�_�e�8�<���~|k���
���4�M�9�Z�U����٧m4�!����������:{�`|Ny�U��'��C0YS&����DY�oL)>�R���;AB�&����Gv
ٍ�.�L���Fj	��� �e��Dc�o8�7/ҥ���0P�U}���۹�ا�׫:W7?wX��@�K��;qB$�ڜ������Вk�[1ܱX:_��G�E��]NFP�:��%QU�3��'_�Y�L�����?��oI8!7��[���͏v
�_:os�Q@�rNMg]+�/�I���4�4�v<�˲�/����Ѭ�.(���&��1�B�\�t�)Jc}q� �o4Og_�y��Mc�KG���s΋�5�g���1�5��Gb٧�׽}q$M+Ң.��'��憎<���z��V�ץ~�8S S�y��1?�M�n�?e��W�BQ�D�����m�z��a�pI���W�L��zM���~9���9+�tM\��LR�t��>5ڟ�돀���|����lB��*^�5^(�_��`I�h$Ma ����>Ƣ�ddq��u��:[��A�? �·�Lq�KmQ
�;�u���W�`�����C^7�\f�FC���JA,K�r^���E&�/ʖ]���'����]��R�(�eQ�>Xn6��g����M�Ұ A�'�}���H�!e-�img.,!\���5T���Kw֜6I�};��{�Zƹ����/$>sP׾싋�WޥT>̷Qtk.4��b�,yt�&݃�H�Wb9���M}�`�TН�5z�Ks�wȍ�fF:i}@i��Lyv�J2oP,��|�x\h�v�c�b����td!ゞl�.gu"��� ��͎�؏��N��l$��
fƸ
�G�p��PoL�f�L�'����}Z0�9�i�S��	u9��5�����\�w9;���z��p����DY���t�\<'����y�z�n
7^�ID �Db;\�ȶ�����@/��3�$�*:mj�Q)F6М�t��"��KW��k��G�4�I��B=��0�R�f-���4'��(Nu���F���+�cL�V��+ʂ��Y��%���o���1�]�b�az�7 �19�[�'�|pω��m]�ب�z�^��X�1�]�NK������f�\a[۫��
��|%>��q�O?�$.C�U���|Mïe��J����˷%�!��Y�|�A��[�h�6v��B���(��*�
t��IZ%�vQ�[��w3����G�k��*���f�����@>�/�_%�E��0R�|��,��m��0��>�4�)�� I�x)��h����*�����4����Xә�W�V?��m�������'̛�קJ��0d��^�d1���5�i*��D�
5[Hf�դ�>��H��)]3 �7�e�m�G(�p[��,��/��RyV�~
�F�dMW`:���p(�fC�&M�ޟ��ώ�ʽ�d�
�v̯De̓���6[�Ӄd�� �k'��T+��ؗ0'2ԋ���&�蚤,ָ�V>8�ex@Y)�^O�Q"ޘ��!:̇Jk�1]L��O�6�P���WM��k��JI�ݹ6�ђpu�@�$f��b�j?+ɸ���r3�"��I=/���)������t�k:X�`�pL��K�%���`��6E�$jj��p��%w�}|qn��'G=3e�h�*Ak�q&�e
�j����-KP��B����<���9Ȃ6�~G�������xЌ�bk��A���  ~�'R��c�����
�08��r�l�4u�<�7��.���N�J4���0N�Ip,��u����g��tD�h~�w�5��O�	p`��b�8��4��F��k�۾>��W�<0>ϑ����!N�&�f'���S������z��]|~�u�zS�Av@�I�Mz������`z�D�Pu�g��|�����������W�ҟȊ.��Ћ�x���Cg�ϗ�Ĩ���L�|��}�����<c��vite��I���iy�Gc��7�] ��J�M�rWK�g�p<f�J�w)�^�JY�����Z���V������XF2��D)�O@-P!����}����Ù$�6C�YЭ��c��T��6���F�T$�M]�z_�nL�`�A3�U  + �f�U�x�'DHh��D@婨�g"�[PL��'�[�Ne��ҍ7I��@R��2f��w��%�#Y�A���ezR�8 ��JZ����n�ǽ�����f����)��b{EB���h�y�u��I�>�Й�Z-��%�v���-������B�k`�M#��\"F�"On\��I/�<d@��)>��ϻ�yʆE�Ꝥ�>Z��$�Uӂ,R��%M�jȨ�R��, �rRd�D&����y�@���Įe���s6���o���g���x��B�W6i&��I�Ā�A5�~   - ���u�x+ŢPDX�"@�%��~���UP|낧=p��qΥ�_D3�6�ik���hdJ�ޑE��B'���ϗ�i8�D�h��v�<������[�:M�_��w���o�P�(�0�{���B��P�*=��֐#h���a�j��Ýl?�����~����Ac���:�"�b�21��w����9�D7��TTͽ�.���l�i�%I����x���nnw�#�K��Lj����݀aTJ���#7�hFl)В3����<7o�駿xe�pҕ���}��N������ڰɌ��I�n��@ԁ�    � ��-����X�	&9C�8��᜼���9e���G�g+�d	��Ĉ�T�G���L�4���`0?�"c<���H��>�t���́*��v��j�$���׀�Ѝ�	{�H�];�B�F�Zɑ�	������ɰQq�<�M�H@ի�e�P���h���K
�r�]W/�k	�q�� �O��H�F��M2(�l�0 M)�5�E��)�����՘�!��-KA�D�R�V�h��ދ�ǰ�v�qr;��E�*}k>�i�v�{l+�B�;H�jR��^:��z��_���9N�vȽ��Y�h�9�`��3��I�ٿɕ)��z�sZ\��� ����S8B�@�����kd�H��{o��ʁ/c��2�@0a� j�T�UE   �!���?�,ĉ BTe����2�rwE!p�X��y��~ޮ�X%%��V����P���N�P=#S�kW��I���j�;����_���~��%	fݓ�튖aS��a�d$G
���6m��JA �8� ��P�oic4� ���@ 6i
�Q�����  p!��6�`��$A  �p ,&/0��+��i�롥T
�%s���jq;еVGb�,�.�+�r˰;*x�&m�&jI�N�#8p�MY��;�]�͙��J\5�#,���Q�Y�2/ڦR�B���^��%f�� E��%���[ײC���5c�C�@. �+(�
\j�T����   �!��90U���@�  PՓ�Y#�ӡ�ܡ��H��1�׮AQާ%/C��5�F\Ξ�PV��D�Q@������y��':	u��X�ʥ8D�5@ @@A�b��Y��p$J���C����g�Yi���#�-L	���}U����&Y�If���eD&��U&����  8!��=HA�EC.��XU�  Q(w* ��N�'K����JdW;h(�����Y��=��
B
�I!tp<�%�ֳMT�9B�/�k����F۰nM
��Yf������<��g0���In,�]�0DHȆ# � �  P���G�K��� �pn@��k׼��Ap��2��j��^��J�c����0�I�N���H�f�!UJX�R��j` !��<�   E��I��"5_��s
�8�լ)�%2�M�-քl�Z�z^��;�F�4�0�IlM�Ӟ��v#×[c��F� �1�gJvi�f�U�J5�� ` � [q$~2��ъ�% R��o��0 �YR)�f���F!���`� !���L@���2)v�@@��w�u_��E9�^� �K-Ҧ���	B���J��:�=k��?�3��7qѩ�{��]�B5��r;�Z_�O��S�ҵ-�!iJH�h`V�p3hD  �扴?+�?������N�-CxF��EU&h����ܵ��\�" �!��)��# H�@ � � t�AOl8�pKK�ZJ�w]��s�}j�"��9Ӡ6��aS�^b�%%bt);����3�s�-|�x��܌QUc7j�Pl
^� ��6趹ؠ�q&� � 1 ��u����m��U�tĬy)�-��-��@	�n��T�Z 0  �Í�   	��`����C��A1����(�%����^��E�H&�&;���Y	y��-P1�8|�u>�9+�%��g\$�b��<ʄ5�J���[�,/Z�Wn{��ߧ�Yz���H�X;М;�n"��0s�y(�94٤�l���#��g�l#Ⓠ̭�V����6𜬝Ö���Xڸ���U�4���f�� �d�S�
_
v�J�C2�6s�fK�L�g�q7�!��o�x> �a Uy0�q�\���S��>��r�C^5��h�Vi��iQ��>M�\uv�Yk7�sڎO,UT�P�D���r�y�o;����W��+�F�D<:��Ʋ�{]������Q�p\q|����b��T^��\!���J��IBH+�5�3@k�CEj2"D�ѫ��òU)�VXW�����<����mՙ����@-�<z�ۍߺ��Zk���z�2��:a@B�Ӻ"����˔�7:J�"��	�Ѵ�3����@���+��]����9�Th��?�g;���c��LQy�746�_]~A�R&0�N���g`~�Ǜ��������@�_L:F�������p���U�Ī���£���<�/|�S���13��X�Z���
�=#�1\_������s`��'A�0�M��[���.W��э>U(8���6�mG
�g�:�o>�l�����%E���\���䮵lIrds*�*����O��s��J�a�Q��I���\�w-����C��!	'@3Q�d��8�+G"�|��%���3��4��	�xs+v���R�s7����@Y^�BL�o�Y�/
��e�Z�s���*ȕq���<+%�%Y,��GY6 g	�q�2j$��J�G;�M��p�/ӷB�6G)�����&&�7�UnF�9�a�k��h�Lk��Q�ಚ��C�q,��Xn�&B��w����D�8�DZv�;�}b����$&��h�P�sp +�dN�)�g����f&�O�<�gʾ�.?$5��]l��oz��4q3!�L���`��aؕ��g氨b���jK�jح[w����H�HrF�]: ���/(π�	���7��v�:v��/�:;��*��*oZ�-��^�rV�ϊ�2a��
���TVh"��	X��xb�0����=���"��M��/関������AV�a����]s���[O�� O�J_$t�)�U�� �~H�'�A}؄(���Kk ��V�	"����|JT� �]��Cw��@�lT_U2o�<�ʻ��)"�ĸ��:���f�R�j}�V��q�{@��^���M��G��t4$�3ᮯ}�$�ڝ��p�z]�%n�pN}�؅�q��r�/t����ė6�_��q�֙i��p�����m��������'T{�y&i?}�����[���Q�N'��X {]K4ʆ�Su��i�W�<��l4�on���t�*Wm�$���Nl&Ձ�ysgAVח��5AJn�Yeye�D�����z��P���V��[�{�.�11f���8i�!dM�j�}���Ê@��!j)�t�j���Àyt���^��ry��x(`<O��������]�{�	K{&Vn���k�p���o�TU���rU�Ec�ɉ,Zpd?���i	ߒ;�D�i���d9�>~�D��و����G)Y�,�Ƙ��j]�;ʾyfg����l7�W���X\Ư-�`3�c�c6�_H˘.�6��i��=d�uL���څ�$~�	�x�X��F����t�9(�dG���0����=��On��m�	ہ�|/�ἲ��D�9p���H(�Զ� ��c�����	!��q!9�w9�NBtC�N��N��GAvQ��9����i�VS:�y*�N���gʊ�Ԃ��jg���T�pP��xjw��� ��(�@G6�M�8�T\h�b)#��Ҁ?��Fw��&��Jd�I��pί��A� �O��w��(gj�f���a�}�d��xK4[v5
ʁ{*ێ�}��v�_�9�Us9����]�b���خ\�bE����i�W����q����ڐΌ���v��MN��OƆ����|�oyr��d��5�摷�8����<��ad�l3X~ʡ̭M�R�kH}�9XIj�F���]R}�������O����a�ϝ��@��#���R�G�	Z��S�ϒ�����(�2��=\{�����GX�x��lλ�׬H�ӤYo$���/&AZ.2�4L���i.�Ĩ�O��o��-��u�$��M�fF:O~5&����<�६����H</�*��<�빏݊��!�m�A���8�����]��B�`��r��E��ܮ"<o�[����w�����k
��=L_��t��8$�e�#���)B��s����p%�	&J纀F[萑���I-;!��$t�r���V��t�6�����R�m<V���/To�7�G����٢S�����m��X/y��&�BG�y  ?�B'R��c�hɋ�	
�����z7��wH�_˜��ǮI����;�!��iҊ1�M�����O��X��V�4��a�@���k��k�\bxB���?/L󌛞���Q|��m�]��te��oө#���t%6�Lf�3�w������JF�U��Hv��$�%�0� "$~GZE	BT���E���P�BH��@
O�z_��6�0*Q����?�m<^���7	;�,]�����J��(��wQ"{\�e%��(E�	�H?EW\fl	�@-�a?�$�s��3 
���=����9�7w�nFN��Ш�	5�}��>�DB�@�Ww�� ����;��|#�+I�����2V{jd���7�O��Ǫ(��Q3}w��̑Ojf�+�T�(cw��nFTh����5�i�p"��l� 	_�ԍh�Jz�ҍ��0�������1d�~3Y�+?p�F$�C&����1`{�����G�Ǵ�b`�x�fj�������J��ɀ�j�z��z�,<�ci�%)�%�*�s�[����Q�:�W�#G����@#A`��Ɛ ���0�u� �AR�%  J ��U�}�&4X�"����R�&hҥW�E�|I��=N�T��v�ǛB) ��C��%��I���
����)s����P�A�`bb��p_L�B��<�������v��
��s@+�q`��T �J�LvP�}�~���(�1��%���	Xꨞ���yT� ,U���p�](\�-�+�~����7p�U���
�?�"~�ddY��?�)$�p���eTǎ.sD�/Ⱦa:*���g���N�| �XC���3�o�n ��g�-GP3�ʈ�GYJ~g0����v�\�DHt8s�e?�gel ��*֘��v�o�D�@1N�K[�c���;R�Ao�O   g �&�u�~1H"LX��@���d�Io��3w�D��mp�mr`hFl��{�lop���0�����xۜ�1�&s?m��PG�d6.���[��Y:h�*3���;����w���1%�É�qڈ�3�Y��}˹sU����0���m�A'���wv�S��j��IJ�I�3��|އѴ{c�Ṽ<�p�o�mz.	���H�DF�~�u���4��eF�>���.\r�mp9�u��|�1+�����5Y�
:��6k��~ Q߈2�7�y'��Ɏ�1֒��gr�-��A�zK�����L\@mq."c�ek�;_����0dA�}N U�3Q�"�&�Y�]@y�aq�,�AE��   = �b-������#Ǌ"堹Vގ��ڣf�$oo�����Z�5�
5�jKn���m@�&�QE��Hɷhoz�F��H�X���~�+�;Oc8r1n��4�)��������N3�b��!��Yn�u5QOzO����c�!ڵ�;ݢn�OLֺD�������p�q�)�Ǎ7�j|G��0�ѣ_��v�B>��ř8�\°>��rH�Ҳ��j��x�����/���7f�K���
轅7�6",���4���r�j�J.\eM0#2��_w��쇒�� ���]'hy��-��N1��C]t�oP�C��)�P�EE�	��������!��50!FK閆hX �+�HO��WL%�>��I&�bI��~5lEZ(�y��s�ɂ���,�k��3s�)��l�v�j�LǕ��d��w�(����
��&UUI��m���8F�� @GV��;�͝⓹�Ұ�e���0.]+�F�1&�!uI��V�@@ !��4�#Sk�,VA �ǲi���`