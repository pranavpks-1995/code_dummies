package nco;
	module program (Empty);
	endmodule
endpackage