0+#�k�����:>���27Y�Є��8�;W �'=n�]�J�zP�*ҕ�l�G)�cx׃����o�ޗD�^�7_,�,�F��LA���Q" qs|7+��X8�[P�`ڂ]7�+A�V�Z�Z��b���z|�҉&�,���v/�E�9r~B6��g�����ӫ��,�G�13/�[(�a⽍YF�ւ��U"�e�����p�^���e�ג�?�2+�-6_��n��K��U�S��*:@}���4�=������]_<�^Kyĳ�I/.��X�Ƈ������h8}?�95
���#G�~��T�%�6�{ �3H��*5���n��ۖ��tD��[o�M%�����o0M�gr]\���u�Z�,~�Ļ�4V(R"mrȍ�,�rt�Q��~�Z���q��~�oo*�9��=_�6	Q}^�\�!�mй$?������9�𹸂���O�hD����\�1p~+�������;	E�#4�lgr�����KM#��=w}�$�u�6�U��ى��DL���z�R=V�t�
�vj���/�R���X4���Nd{��o��5C��Q��>�<�N�o�QS���,��%�Y&��Z��Qfܥ�G���E(��8���E�a ��QQ��]C�Z�O�Y�#h��]�W�5���LkJH9M�[V]׷�~��	uܛ���}RuÍy�\ك�:A���wM���YD��>��F�X��2G��}�h	"N�"�HHK�� )؂(�X������s�O?�u����-���k�^N�Y��oy���_-�ֳ p�><?Ȯh-�!I���5�3�WJ2�|f��=,	�#�����t�|��cLk�����%�ǭ�ATpM˪P$T����n��>C��G��
�Ղ�ԑ�9ZGZe�QQ���� ��"���y�a�7/c�RB�.V�="��M�p�ջ�i���7���&�x�텗~��E��ƳlP��P�(������Ŷ�X��
�U�𿥎���g��W{!N�������W�<��M���]�hT/��~�4�/R��yR�b;�q1(v�hўf�[�q�UhP�3�P��#�A?n<'w�ҙ��C�߂�i�����֞�����_1�؇��2QU�56U��}$V��&a��z�����3��6]�A���BVKt'�2�۞V��x���}}��o{o����o7=L�C����=�ie+��Ȗ���oK�ok������/�B�����<�,L
�7|���ћX��M�J�ۙ�nv����1�������z�E�M�Uǚ�`D[V�L���o0d���~s�Os�rR㻌�cA�����V�H�S{nyo�ZP���o����v����<y N�𮟏j�J���	tT	=w6��Þ@�	`�<w׮�c�ݷ���=�9n��@�nR9���W�
��`���\s5k�} P؃e�1�bǶO �����w��Eo�$͟��Y=Q1A�M��>=Gl�Z=�r�r͐����,���.�\zk�ge���{�{ώq:Mwl^�>�ۗ�G���t>vA���6�lS�"��ŴHR�����q�\�;��[Z;[i��c~@UR�k�TG,���Oޑ�q-�|
�Ő�XfY��P�&�3�uZ��h�6H���a�p�����p��U�מ[~7{`1�T[�	ܬ8C=��������-T����z3�ƽ
���8�Hji���rX�ⱳ����#�>Q�K��6d�l�Cr��.���_�A{���{U���WDf!w�'�+K��N����g)��WP���(\d9s��)�A����z�Q~-�ʒ$�kH��V}��T&Hш:ں1���~�,=%k>Q�vA܃w,(����L+73tЉ��\���
�қ�Q�7�bf����7#�:CH-ޏU��D6g<+*����.���=(�����J��ʏ�Y���?��_ ��^�<~}[��a#zi�ݬZZ��"p~}�]�4�u��+o�@��j�5���ۗrQO�Z�Bh�Kw-@��\:|�����pR.�G�,\�+��H#�zbvV0,�뾱&j��%�B.L���%����(����pߙնA���I�_�h���Cr�2�T�:���u��$�aW��C�*�xK�t�Cx����)́�6�ꇢ0;����S��i墓*u�3l�{��#�9�3��}{C[B^u���7f��%�K�IM��P���	]��j��3�������B�ښ�N��;y��o���ز��=G�l��H��ctS�n�Z)���99�A�e���c`|D�H����9��jz��=�e�Kщ5	.�E�d���Y%)�6[P �Z��r����h��I�!IO�	���S&�s��� ���Q.��*P�84�֛ �� Fx�<!�d^)B�P����#B|Y�@{��SKS_��?��fGp����ž���$>�����.p������\Z��
�<�+�`xrr�O�[C�V�\}�&�T=��tnx�2����mt�P�(�6�e���q݀��)�#:���i|�QV�g�o>$$�����f���M�;�k:���fFF�@�Fh�>��w<$�LK#�`�8��~��
��\����7.w��#��~�B�\�v9�@`;D���zE��-y۔�nA��fv��IAht�Nˈ� �n@�N��v��8!p��ȫ8��Ʌ�G_�srI�9�*~�S��@���65
c�b�����4q� ���z�7%˒]B����{��F���m�$�J�mar33A�@~����rKƕ���jw�N؂P��]�ㅋh}۰}����|��+��j���>]�mƤ��	9���f>i��}O4�B�G���Sv�a{���`��J�������D����n��bv^��[8�ӛW%3�K�Qʕ��է�@���ddv����87^9�pĊ/��K2MD-��mu�Ji��#�8��)W�;��y�ƥW����cX~�� ����gg	�͑��x
&k��n���P�|�1Ƅ�DH~}�^��{��ѫ�ő�#;�r[�B���
zQ�;43�5����9 A��T��(�T䅠��1��(Ma8[R$X��(
�P�W���s^w�NRwcm�K�T���1�ҒW��Y���.��p��.1��0�I��b;���:�s썬�ƺ�l���Dr��&֤<Mi��9�I�t^��q{⮿� �����OGC̊C�#�[�	�t�eQQ[���;�������x����o�,�b>/�dv�y"����|��t��,)l��?��%���YMc� �z��)�m����F>�L|��ݵ���1;=�kK3��`P�D�_���|Q��	5�����ș���fRK�ߢ�u��+⧢>X} ����'�=�փR�h��0F��vGυ�rM_�47�Z��v��5�s��uޫnHr�>��{��<BߦV��D��*�A�o�������@7�w���c=��q���wsNv|D����>/����U�4e�[�JMJ ���Ld�l엸���v *��������rwSW�~�#|_T>*�oP�/��#2Y�ѥ����`_E�̣c�"2�6�Вh�XJ���15+4"�![!l��hN�=Y1�fr��ŀ�lKM�T�<�ftc�y��[^4ݶ�=��i���bQ7���9t����wR�`�k���"�{�F�,E�<����z9��<� &ߘZl���Qp=�"�,`��J��|u��z[�:��ךS��MuB�*��*l��k��y0J�&�۩�q�{� ����@,l�T?dH�F�w�`�A�=Ԇ`�E�7p#&k�K��L�xB��.����ωN��K������2�8򐂱��%0�G+R9d��/qB�������ٝ�;�4�$=T�8]±��h�*+��|Z��)r=5=�+�؎�sr����1�^��~}B�R���ж���?�����QHC�u^fP����c���$WƄ c�%���!�J��d;�k��8��}zTF�J�A�L7�P;�ƌ��T@4�!���&�ZQtxtS�� ��DX�Ӛ����^�]%���嵬�
�<�$�<�#��)���Z
�~����y`�F��r�5nT�A���J`:h�����\p�!C>�0.I��lt ��N�fӋ��8=D�6������p����o ���,�s��dK$�V�}F=f���;{��p(f�Ӟ���:J��Y���i��0ێ�	�����2hN��jW�n~B�Ղ��!Mf��-�栀�-O���VJ��QV��[ �h2��>���˳�p	��	�M�M`���B�ܵ�f�kl�5PW���4����x����ŌD[m�%,r�*$^�zi���4]����x�F�D����h�����m[ʲ*�ٓ�^@�(�������h�'/�lUm�A��O��	��]�w|�;=��9<��_"3�A�>�7�lY���~V�31a��1wMŁ?�zfY��K!���� H�GũB�%Z%ʤ��E�3Px>���X�fN��L�F��L�@���N�O���e�:,������!���'ٽ;Sn�q��s6ϝ+� Z+c@X����������eݺ�~����7�OQ&K�{v��������𝺻�G���"_s	qT�*��|�)�	'�:�Ve�i*!H��[�$��Gu�:W{hsT�Ͽi��3��(I�J	0�R!���JBl�\�����Ucq�oRn�P��{�4:�G4�c�NO��l:tg,a�#���˩G�*6\~Fѫ�V��ZK#��[��r�^J��eY��˨tb��湼����n�G,p�Z|�<�N!�8b%��؜�S�9H����ޕ~��SIb�7+Gl��	$fo	W�d�~>�`�� �
T=��Lu���:oˮ�a�ɲ�p�>+-1�o�U��<N�� v���wC�������Q�&�z;?[�|$Nn����m�����J�VTf_�X�Z�)���Hp&�]%�!��N�kV�t�]�`�O�q�c%.VҠ 
��+��?2�zcM��>�ә�LJ�ٗ!K:�u�?���(/9�o�4{�y=���2��7�B�q%�Z"Է?�7qBK�3.[��V~X���m��d�x��;6�8�e��6�w���[B:�A�Zz��U���7���D�o!�
,�4�u��k:�� E�R�x�����x ���*�.uԊq5d靧~�V:��,@�09�A� ��Y*�`&�V~N��A�ֲ��%n-���rb��;Q�%b���vXe|u�F��5.���i�������-E�����N�����Ά�&|�11��7Y�\T~�l:��EU�_�@�`�k���8�WT���C����&�<b�v��u�bro�*[�������My�|�����C��O�쀗>��ﯢ�������C�jx~�]^�{{�Bwn����j��~�M�iX��	�}|�Ϯ�HY�P�Y��KKsK�X6�sV�]�0�,�K�Zm�K�܈��>���[��څXb���)��A"��a	�d�Q�(^7=b�XK0˻�B�u��J��Q  
���'RW�c��͆��	���l���JM�Z)"��os}w�1,}���i²im��������	nS,} �;��������r�Cc��\A'J�x*�2y�Њ����p%��.��z����F+\��D��u
.��ZR
�D_���6��� ��[��u(yq�;ұ<�YYi(������}��B�d��1�w����.���p�������hBbI��c<�	r��f��Is?[��m�i�P���M��G=�ؓFs�	�\��%{�ʕO0��}�0s~o`�&�Kf+=][/�P�TRr�6Ԝ�~�B�������FW�1�aH$u�8�lz��'4|��g�`���(�N�˒!���S�F�}so a�{0ٕ̰����rF&�f��8�0s~ *��������<sГR����T�~X�F�$��}R��@i�{�p�߫��-rఀ���e0_RU�<�R����Zu���]�^�Ic����?��9x�9�9��^�7����q��*��8��@�Q?�GT+��
��ψ>j��#U$ȓ���1�e��h�0��`6�\h0�*ױYK@�����9�� ��̖��_�?�/x��^L}�+ķQ����AGϷvc���/M���i1�GO[n�h������&�養D���vyO�C�@R"-̣�SԪQ�a�-Q\\AC��]�ņ��[O�� ���z9�q�\8 =V>����$����4��<	�x��Փ]V�t���}{9A���_�9i���(���*sY�f�����z�XqQ�����qű6�N�7��:m#��>y�ߵ�"���O�MC{Wx�i��P�*��x�w��8�ZE;�R")�uJ�|^ְ:��6�bU������\�N�ʹ��� �\��ra�&�Azyh����A�Pg�~��OE��s ��,�3�����S��<o�w��8���ۣ�ê;�j�~a(a$8�p�^���73�hb�[�a��z��J�xU;���{*�3(��f��ߊ�+֢�3����UV�܋�9xR�f�#?�P"�Ѩ{�ަ�%.9�Og��!�B6Q�9U�4'��}� �-ZPQ�Q�u
��v/�ME�?��J�]� ��
���Ћ58t�糧�)5�Y},�ѲTk�UH2��b;����Dz�q>�Ͳ����e2�	/!!ּJ�f3ギ��>�!8vXj�{��!j����F�X�4�h?�������"��X�v�=y
⋯�.6�~�
�$��N.���yZS���$y�H�~�l�4�6���?�n�kd��%�@����,�CƵ	�}/��x�C��R��p� {z��#oN�4?��=�m~��@O!C8�j휾ς�T��ulU�	Y	?�Q�qoT��G����4��%;�t�0����ziL�+x���ꐼ�p6=�]1���j:Q��J��٥Z������]>/�=�N���ƊZ���E���
=s���f;Ьz������ފL7s��)�����d�;����Ի�T��=����i�(��m��G=	�٧*9�<�y�"+v
�+B��NK119�:F�h����!��p��?�f�b;w��F[��>�m�'$�"
�+��\6����� :�Ny�}t��n�$u�q�=yw�)�9�~\��=�pX�����@�E"��A飘B��(�eA���j�"��z�$L#�_�.U�g�p#�E�p4�S���-ŧ�����"����7<�L�БJx�u�]�6��y���:����7mm1��Ñkg�|�,j�L���%���}�Qc��{�c
{mv�g�����R�� z�J�Qn��:p�ĝ���Hr >A;���mX����W�{|J ���T���M��������,�@�`v��s�B�-�3��|���咺�<����ɥ�]}��W�*LU���t��#���̉��qދ��,�H������ܫr�f�̔%���՜D�cϷ�.]�0�]<�����){UV�χy.��V����.!�r�?oo�T
�;���p�īD(R���5�ڎ���J�mJ��@�6H�Hv~M"����V��W����W��J���4i���Z�&R&Vm,���b羃0������_p��f5�p`�̦p�w���d��G.�Z�
L�Y�kYV�ʷ�nǽj]����aW�t��.gqmU��0�[�m�x&}T���X�m����c4�VT�C�B�g`Q�>�J���7����rs��v�RTT0���gq�CJJ���!�7Q�A��Y1Df�#����ys	`��?���~�8����wC�ޗ�&"6��
�.,��@Q�j߯���=��^��Z�"����뽌~:�sl�buLe2�;��<�>�b^�.���)������Җ�]�) ���
��3���¡��� ǘ�T�P/nm��c0:�w������H��)أ���D_S'�+�*�t����՘���:&��c��n	D#�1�����	�n�G������au����V�AsJ�� M�Ys��j�͕��Tq1���6�H����e|����hX���!�[v��jLG<7�g�B傿�✿/�7^�E	9�t�B��Ǐ�`/�<�Ua��ҁ��Љ��R�L�6�9�n���J�V$YOz����� �y�R6^~� ��T��Z�rǝ���k5D��]X(��(#��Hׁ�  � �f�U�$�Y(�R�v3�eo�@��I;,r����_�]���g��F�=�H���C�v��Y?���Vi�Z���G���P�E�]��>W�0m\{w�����MD���[5���������-a��VS�kc@o��>�}�B��L7Hj|N2�mF���Th�f��˿_-��z�B���'u��0ℴ���Q�?j����>�p8N�%U��o}�"#AP(NR\�����\������^=9��Kr(w��0@X�:��)`nA����w���k;�Q%���w�0�����5���ϔ�����́��'�'�jZ�)��j��i@���X���Ѓ{�/��Î$�C��ʔWj~���É���u�^�_�Uy{��a��`�#3�+\���5�wL#��lS�-�{`�K����?-
\�1h�6�&�ul`�z�[�)ǎP
�6��0V?���;�V0mi���0����F�o���;p����JI[5�~��Z��dHu�K?؜$'\���V:��j
{�@^�IW9K,]��4�+�;���i-׉�4���p��9���}�]�0Io���<���&),����רA�|�]�;mQ���?R�%��3��h]���,�׺��Zo
e�qM���j�*�@;S-�ȼe}k�д��̠W85u.���I�q�0jɌ��F��o@�s?lJs��$D���A�Iw�_#፼�ǎٛ>����`�+c������Ēi��<�F�2��A� �Բ,6ͽ�ͭ�yc�<xotb?LL׌���w'&�Td��dE���0����h�9-���`0#5Jƥ	iQ�ßL�ӳ<����JOB��x=���޲�TS�-�<#�)m�Kj�>7{�:y���TN��@1/vg��8y|�ةt���2�=D�����نBI<�Z;{&��X��{�9�(G>��Jw�
r�|���U��gl��B%y�ٚd��z���b�M"�@m�zU\p��L�Z6��Y,�I�AHJF?L���5�y��E���|��P
�'a�{����R� ���b���F��Sќh�3�d��y���Jqz��X�#�dŭ�f��l�U� }̔%�����*�Ög�O�xKl��NQ(e��~�l�d��iDI�5��!�:2�b_��!o��6?���A����A��]�5kט1�uA�r���i]��w��	?��n������ԩ�L���L�1]�u�*o�U}��ܣŬr^���Y�����$�-���
t��6%�C0���ݸ�G�����.�Xo��1+ų�r����?Y��C�����9�����^5�I�陷oV/m����@���3��D�'@�* ʹ�GjP^��I��������̗=�0� �D�ǫc���[��2�8|EbM��U�h���ŧ��T���:�3�	�;�'��f�y�٫7�(u��W�3�B�q $���0����É�)Y�@��Sx���]�M8{\ʰ�ޒ�M5���T� ���V�j.R�?/E�֘���\L����.���Aѝ?�($������[b���cz�Ұ_��L�{0�Xm�8�Wu�fI6��Y�\�P91^,����4��(īX/�wy��cp���b�b��Ea��{��$2P���&���r-�zʲ޾ś�3�]�5~��_|��@ޭ�>�|���>u���Zb�~� _Ӑ^=���.�"����!\���#f%qJ�ҝ�D��<��]�[F����]5����}� ^P�Q���l�G��Uc?`V�x�J����=���u��
Z��zMJ�y�E.��q�?)	=O�.<)i:���y�}�z�J���G[$524dK���@%;��HS>��hc�k��F0!i��`Vs.��0����R`=V�/��IKBiQWk�[�P@�=hձZ�#�ƈB8h�$�I%��T?8znߙU#�Z��=�J] %�r@\�G\��Z3�F/����)�w]��@Nd����,�{��>4 �(ׂ�.�;ve�M�������\C�l���*<��a�ω�S�F�SmG��6�Ń�*�[A!_��N��c=�sv�\!7]=���x�j��1��Aݲ�&�KV7�I~�[e/��	�ۊZ^�{���M�\�X4�����B}el����x�G�.��-�.VOF�L�g�2uO`2��P�2:��}x�Ão�,��0r!(��eӚ�,��P�Z��iinD/%+N4!)��HC�'   ; ���u�$�d(�Ы&+������u��8Ag�Q��c�+E�Dng�f}�и0b�1܀q�!v��($�E�2F���������s���g~������MSz	���{�0cՌ6:s��Q�"�"᠍Ĩ�08M�l�t����>J~�ʏ���et5�3���c-��~&���V�iA�|=g�*�'�otЬEKsT�l��4�ϭ���⒖�����Vg�j�� :��?�l��jp�*%�H!������m�?�1���i඀�p��*u;�\{�&酣�N~_����0����]b{Jg|+����As	#���7��:�X�Ş[I�޳&�"�?���@�%u��Ȉ�?�X���