���*g#ꀡ 	Ɇ׬�����_�{[1�-�����{�����m�Q�Wk�Zc*�y��m�d�~�L����5���9��-�h�q^ET�KwYu��f)��TU�2���s^�I@ �҅���݆��8��Bo�P��'z�O���̿�z#����}9��z���f%�-Qn�K����!j)��Ù��j G��?�y(X��<<�'f�Ղ����> �� �_��u��G��w`N��I��"�_p���� o��T-�X���A=ŔG��+?s���������&,*�?���(��K��RUcxp������)����Kc5�k�����<���d�1�2�Vy�ڧ�0�
l�<��ڵ��*T���A
C�����`��j�a�b�>o]�l�N��9��pJ�j b����ls�����N
?��(g�i��uJ������[;����!��(��,�?�N�H���DO�{�����6E��ݡ�ԏ��jӔP::ZhC��l����E��g�y\9��e�mI���ŕ�a�X:�1��b�׳x}Iy�0'�|+WU���5���u����K4�㣴m g𮵋u��u����2TDT&�"#��t�k��.`�IR��;�&����E�Ɇ��/E�/F��� ڕ(o����9>f�gf�"�,���.������MX��gS��*��r�#��do6�fC���A�3�sr�*6F�8'F�h�Yc.���[��,7%w���^�Ա��pq	�m��Иc+�V���&U3tH,����ݡ*����{u�#�ԉ������;@H����{^�4��)tS��m���6Bj×)|qy{�o]�D��V]��S��O�̮��4�Sh�4��y�� ������?%h8�Y;�n��^z<>���&o8Sb��x�����ઝ��x�M�_��"��wa�j����f�۳hU��`?Q�Dŝ.z�a:���.\�����\J%��>Hh�k��m�T$н"擽��xH
��q�y���R@5�!�*�G%����975���
�,'���VA�D�R����_��Qx�~�u؍�4x|H�>Y����P�O6�6�a.���Y�� �_
��Yoٴ��`����GN{��8����""������`��XJ0�D?�$��6��p��� p�:���}_=�1��K!؍�ם�E�GQ��4�K�獛�a�.�a5�O�vc;k�,B	,�uy^32�L�J+�4��w]xaS��V��r�X�Uޕz{:t�3�6�j� T��H�̈́O�V�;v�p��QȐ�>������?���������.�+p���4��y
!ɱ�C},�Y ���v�(��գl�'M&w0 �<2��-�i��S&�����&��h:�{W�eX���4��7|���"~�oFf������lD��^@�	�c�-<�m�� ��{n���U.y���ޯ�z=�|���R=���l���T�ji��ew��'��}��?h4���P��)�6��1m���K�$�9Y#��9Z�&2�)�'T�l��R�\bX H�����Rte���:=,�n��dy��~��G �8׳�z��Pe�m�Q�66��F��e|c�hn6ܲwg��9������"r���^3�5|׭�$��F��F����T�{m�b�WϺ'�1��&�7�5��dw���`P�_R=����G���Ek5sy��tȱ��갌孆����
Q/�4�1�v�?���eP�����196��t�o�L��G30m(Eo ޥ�g�ii^I�{����^��"�wc��◀O;�|W�������y��E���D�y�4mQ+FX��Zw����:�lF(旐�`��}�.e'dq-&t���_���ǹr4aҏ��v�)�׋b�vR]q���]� z;�a�[)`E��#���	����m)��M�ϡRF��!=p���T�nMnʶR;����,h��̘&����`�5Lf�R��͚���uV���e���q�&�*��9��>M�Y���뗅�U�C�9�)f2�	�n���A)J	��0�}�T��ԕ#�6{iĽz�U�uA�z�fi���ưD�U�
E5��!T��P^W���g;;`U�J�9n�/�g�$�V�"j�vb��sb�l��ryZ�����1
y�%��^cU@�շE��_&̈́��D�e���)���8�#�g�Li��l����N_A�Dӟ��l�/�hglG�b"�KJ��0q/ܼ/g]ȳs������Ϫb%x�@uLt��w�zi������1����a�\{�f��M@�x���-��e��� �ò,���K���m��B [/�=(��	�\.!��PÒW��m1k�g����q"�G�kl�EH�k  @ �����,t`�����*YZ�p�6]���
��17�O��!�"b�@�(���ܚE�oGb\�c�&z=��R1@�U��̬D�f~�a���dweZB�z**y-�b���^"�a��#r*!Y��l$���c-�~�BI�,�k�[L��?����0����������oA�-��njc�z�����6�$���q�l�H�#�.�WC`�ú�C���X�ʿt6ޯˌ1O�l@� ���O�>!_���h���x������5M5����)���ɯ1Eܞa��cN�lĤ�B[�h���K���u^�ORB@���K����mFλ�o�ǣ�L�F[ȀH�\�4��D0�^[�<I�"�	^r�7(,`y2W7q�X�1N-Zqc�k����|��h�ͦ.9QD��Ѷ#��e|���/ �����O7�9zb�%�/������&f+��殺["Ď��;@py�N'�w�HV�!P�dfQ�x#��F7�+֞L����~ ��-�
������N���`v.�	o�����LE����c���1����99������A�Յ�<�2�U*J���.��x:��a��&�*�0�nJ�#���%xE�Ê�!h�=��M������@Ə��}�!�mA�����%`�$�@�*w��v���pn3a��mݑ���d�󤥩���~����ja�к�.�ʡ�.�lpT%��j�,����ˀ�e�病+��e����K:�}��h�+��G8#
�|��ičT��U	Y���ݮ6��m�;�ɋZ
�Ȝ	ׂK:Ũs���{���݄���\ՃͲ�>�/� m�7o���Zk��_��2`�5ء�hIL��v���"�A"<�_�{ד��Tfk����q[k���~�Cn��X03!�z��̮Pg=:kDoR�ߵw���e�s%*{0�c��߽��Ӷi�+�$yE�w�}*r����O	*��@]
�0h�9��Ḅ`� X�+�xFX���eiw��/uFv[;�z}���k}5$�W^��*p��l�G:/�A��/�j���pr	Oyn|���Y�� ��W2��<v�>C	+50!хo��k�I,���>��Y݆.�].<"��ېrC.wL�V�.��I���H�ekOdo�[�)�x�?���Nc��ɰ����2�M*5�D��?�"�K���n7`�NY�#t����� �ֱȮ��� ���- �~!��7t4<+������ӄk�3�q����ێ��W��A�˯�u'͵���`@�Q]�����M��2���\.L�4�+��K��/N  ;�}���x��D��    ��-W���U���&y,�!��/"���6�˘��6Y[��[�dҺ1�Ҫ|)��%�|��0��4�j�Y'�m�K$������?�2f�iP�>�W�-#���Y�x\wUۊ[ý���;D+��$Um���h(3d�X�V�Lq��^j�K�\ā�!���S��!��t���ރYkD��f���������#ϥ�e1�'2��4O�Ru�$�<���oA�v�d�D ��"��gIl�K��q/�H���O3�R�z�K��֯i�èQL�XXN�&�tX�I�[��R�n��.х�K����"n��Y�������zT�Xb���Y��^��ڸ!�w)��!q$ �7���"�<��82i��0洆�E4!f�j`��`�צ�f�1��)��T��k��h+������Y�^��7�ח��l�Q��C(�9�#��s�bBd�r`��|��:f+��-�=zq�(�_h�t�0����*É�^23�94�)@{ l�4sPʈ`j-t2��n�|\q�lUQ��Ƀ��G-��6�`�5!��2G)9��a��߈[�)U1r�wC$�����NQ��
�I*�{�õ�ª^;á��tsYf�3lT���Z��
�d������׆Z!���x��=�1J��L����6�]�� ��0)9!�+���2J]��wK[}# ٫�H��:�E6B
�����S�͏�ؠ(P��j�0d�,y��{P���N��!��v'�)���ӆ�BF�0t������S��b�xDIc��k�T�2�4���&P��/3��%���k)F�k�ι�Z���gisK�iy6���>�5}J�g<Lj=QR�R`�������3���G1Z*S��j;h$"c�'��?sȑ�]�0а]��e[�`M�>��~�7�R���t}�_�K��J������cԨ�<FX�n>-b8��a��	-��Yg��s�.�\n�7np�:}@�'�K]��U/�E�D|d֚��j��>�B5�]�*+��H�Ĉs0�EN�	��������!��EL�"HZf�  X��H{�țҁ���C3�Q��qvKT�]��)M��%1UU��	l)���uZ�ə�Zzi^:BiT��+��Þwn�fG��;����鯢�"��%Y &�!��  �\5�	(�h��{P�� �] ��(YD���49 iFD�Qk�T�"TrP   �!��<��"�R&�@�V,� ������"*r����R�"L��6���0AS҇2k���O�<Ka����UD 'pj�5�E�)��hX����n�
��]�ɸ�5���`�?��-Nh���T�w�o���`����	G P���P$cCgO�9~��p(h�:�W��o8 ���HUR�*�  !��$�+ �V� ����@��|%�'?�<ψ:fT��:���t��d"V΃,��h�S�L[L6�&��QP3�2*�l^���&c�c�%�c0 �A %�X�ך��u�\?��߼�����'x~�^�P	�%g��F;���C^������%A  !���L6 �)�(����%��μ��V$���' )Sut"smgfw̎(��1�\Ƃێa<r��j'�FH[�T$
�.I� �Pa^�Z�%��0@