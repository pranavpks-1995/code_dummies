�\~�z���-�1��
c؋\��wH}{�����'�o�t�������jռ8��˖��-X+M �h�*��Ѻ�ή;NJ���Z����{�E�a,�?|^�g% ����)�d��M�|^͞�|���Z)�2   !�h�UW�C��k�ԦIob�K�)�n��c6���;L��jE&e;@���A݉��X1���v�Q@�DGh5n{��$����1
�M_I�����������-���C�:u�H�͔���[.�n��з��H����>8,�):�g�.�V�iz~r*M�Q:I�va��T�)h�6}Gݤ��d��|�'�T5���5֑�9�.�	BvL-!�6�J�ˮ�mW#í-���� -���J���I�ꈾQ�v�Y�5�(&�xAU�Z!��gA�s�Eu�����lh����i��\Xh��ԕ
��q�ꑯ#��,��Qae|_ ���X�$���?_Rd���Luc�;I�	���!���C`YdX���Ǆ�����(�#�!{y2r�S���F�^���-����qDf������;7���}g��pPL��1��"ð����A���|#9��E��A���i��d$�F�J �lP�x�� �Qݐ��p1�H��#�Q�_+��Ō�{%L��oS�o
3� �M�L!hP^jj��w�
A(~�SBa��h�8�r��=DJV ����\gWe���s��}~��|�3E���v�4@��!��B
_uK�$�u�s�����2~< �Y����Y��ֈ�~"��}���g_
Y�`w�<}H~/ߦ9R�%��)��vd-�Ϗ�
�p赺t�m����F���W��iQ'v��K��D`��գ'����h��-&����u#
c�{r����_���f�NQ�@�Eϫ3_���ѸL7�%��VfYUc�~�{jdF��s���
� �Ӏ��y5�c�p�"�8�-p�
�c����*�&a��b�����X��t����]Fm3h��D�l���ȕ���`�ι��<TI5
6��� Au��NG�T6q����r�A���+�n�o&�+*�!f(���&]�%p�r�'^�"DL����r��!:B�0-�x���n�$���=��+�Yg��u�5��ګ�f��c�=#�l'w6Y��`�s��l� E)���k'g�E�ѡ[����ڊ2�����N�C�ʄê� ��ܾ�4Bg>	��*�M|��ǻg�tw��Y�5�ŧE��M�2�z���KCN0{�2��}�����
�����xuhJ!A9��z׊����������
ۡ�F��wyK_�3>�0�ؖ�yb��m��SG�M���W�����Q���������//��Ӂ���uy�f�;+�ƺXe�i )�f��7<�#	#��/�gJJi�)g�, G(�@tjZuY�ݼ�[gL٨b�����=P�!a�|����7����DPZt�{	��|�Sv��zi,���bzG�v��Z�A�O@m������FA�u��غ��.2����,�B�GIT+���@�:�m*��� �3�r?.�