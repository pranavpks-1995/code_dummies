�����tL�ԧWpz�j��D8?w��ؓs驚PQ0yH,��M,�g>;�%	G�?�1�0�G=�ԑ#�HP�B�4��`	�_�S�'��$<���`'9�xQl	Ȱ�.�������AC".̊OTj���@x��ͩ�h���׌����={�S�Z^p��P�������WSSr���Hw�X!�В?�ӿ��G�ѷ��x�B,u����wТ銝��5�!|�|���Ff��("�t�r��%���C8�����`A9�ʿ���G^��a��ʉ3KD���P�'	�B�^m�51.��*-��]��kR<P�mL��(��gBa��U'�*�\������9	|��z)�w%{��w���Ϲ�m��@B��	i���A���!�i�E�.���>�C��p�%���Z*���mI�����K"��Sᬣ�s��e�[􇠧kW�;g.���7װl�ǿ�8��r~\�����<&h�&�C�e���ꍫd`���#��$�(��}��C���,<�#�ě��w"�K�y�7=�zFd�&�AcJ<����>:�A�}�+}����	�s�Ui�	�o�2�9��	��c��8�D�i�-D+�?�(X��s[,��ђ�4 ���x�f�'�I�I��%WL�R���!*`,�|s#3��v��\%KI+�(<=#َUo_���gc�f�}�Na���U�����ƴ*�Npg�4푇��s��	�ݩ�B(��_S�Ǟ�EA[SA��#��Q`��֐�n���Ux�r�m>7����W���-�Zc��?<�jb�}1ظ�;��ŏ0�7����� �ƞ��G�ۍܣۨ?��-��yNX�#�ZE/���pZ��?Kr?��-�9��TJ7	 u�� ���h�Jϟw�!�di��k�bC�Oa^t\��D�U��5�ǃ2����*����X!\_��n_8��$w�qW:�H^ھ8g-�u�e��\�٤���|ނ����ε��r~��;§������k^^f�h���AɎ�����E����#1�2U������W�}y'6s����ߤ���Z����i/L�j�(P���Ò���/&a��]=IA�@��4.%��7.r%<�Z�6���Cx~�ٻY�|%�1x�f�{-|zS��P����qja��NF�8=,���ְ[�y�ÿ�WdJ��q6��.x����:�PZ�j�0��w���Mo�!�����~Z�5��򿶃���#�;�����"�m�q��Kb��24�a���_Oɷ�y:1�XQ�)��m(K��
�_�v��<
&��?�{$v1�Y4� `I��F�P�[2Pgt+�i��j��-�����Ա`,��W��)>�5�� �y��1=6c\����Y�?�7������ʓ�ʋ�e{����w	]!�������ޱfYdٔ {k,��X�=�|�-Ph��p|@ͮ�t=<k�n[�� 8��LC�YU�'|�G�����8�k���luJ�!�n�G�^�_������ØX�tz�E2���jxٙ�']o5��t���ܡ8_~��/W�HS��)��o8u���ꝬO��ws�6&U_Y .G���.�3���uD^�'��_Ad�iι�.���MvC��YI���b��3g��;���x���l���6�gS�H��>�'1��T��\-0��GhN���M�Z�����"z����3���G��]Esa�~���Ώ�HJ+�� �٤b��T��E��O=���J��O��m;z��r�X_�S�_"�ӧI��wtJc�mnv�7p���/��]
����Kx�,�o��J<[6@Y���aU�Xd����%���gGJm����M�q�nz[��/4�A�J�� �q��0��B��X�Q� ��<{*�y�a f�B8�o09�\!4%�"� �HH�.�RUf㊵/�p�ה���Sy�a�1�D�̇�Z@�v��^N``	����D��~�Ɋ���&ZM�m2�ܹn ������$�6|?�V1���LX9��bnC@��9��A8�k�������EeQ��O����e28��f�	ؙ�[�>5�Gmܽ�n�0�����W�X�=>�c��Jr:Rw��w\n��1�3S�-g��f�lB^�FY�eB���.�3$o�>�����Y	��V��E�K�C���\���1��<�����E|͚I�'��tÝQ@t(;��'V��q�[?W��l�I���$>����p\��ԋ@8"�%����`q�V�c����j��܆露C����x��/����V��4^Ӓ��}�u8 �B�L|���7VZ��u��=�E�7���HO��g-��B��JV�.&�ոuE��0�:�7J��j�����[[��;2P�3�"n38��Z���mՉ$�mKwd�%�m����P��P�'�.M��	��ϸN��7����`o��HWc@��� ڔ�
��˹<�>z�9T�~�gk�u�VG�k�A�r���o�CP��H?`��B�'@�Z�dDQ+�K]}6y�;s�`O,��O����ZpDä�S�'������$'�s�d�1v�:����c ��寝'�2�g�T�	v��������_�����I\�h^^	<C�����<{f��h�N�c��)����W*�Č�YN��EǊ[���6��߽Ges����J��&  
}�%RW�c�M���� �9�P��Ь���Ғ�FGѫ�e�Yr�:��� m���AK�$�v� g�A�|y��U!�n�����8����L�_���&	~�x|�V�{��ߝ�j4ˀ�~\��/�v�٥d`�R�B�������
=q�W�&~>bbg�Ĭ�h9�ɟ3Lc��3��=a�>]�f�������pMU���?�T��Oɵ�O���^�X�@E�(�G0�����Hc���f���_��UY�n�'G��6�p]��7sgx� �o�6��S&U6OϮ��q�fC�8/_���nM�<� �X��y�_Lx�
x��^Ð�ig��dh�)})o���H3۵O��Fn� �Z���9�m�חcQ�8<��}�@gv��9�`�,�hf�h��R�2���]�����Wx`�,;�Q�F��ۑ�ܭT)G�H���s<L���-�X�)3����+�{�zEA`�xPDF�����χ_�b>�а�A]/�Q�7I<F��@/������*8?nFE��:I�ʙh?�"x��� ɨp����D,4�h��Jܧp
�D<=�Ȍ"B�s������.��$��M���?D�Wr;��R����w����+��B_�3�����w�P6��Sǈ@66���@ۀ֚�s��69�c�&&�
{���u��07�zzb��g?���ߥ�_Wl�k�x��mm�+��?��]E.������,UC6͞�E��͓E�6J�b���z�1h yaz�X�%����9ն�u��Da.��콥�v����?O����
D�@��n��Xk
��?W4��k��31)s a��i�1f��������.�V؈B`��6�U[�G�7"[du�>:�Z;\�����}�,��&�Xɒ|E>��!>�<�ITB��y��XG���܃j�>���˽ !<n?6���ٺm�9]ٻF3
GB�YMqj�xez����T`�q�K��ǓYeD=
��C�*L��Ma0����2wU;]��y����9ś�4�Hz��S����Nѻ��_ٝ����qd!+/󵋴�����Cڢ�Z
T�

�é ��3����:2h�KoC@�GY�g�����8J��9��m6N� ��0O�F�G1J��G���K�8x`�����Dw�z�9���^t� �W)��Z�	S�S�~�̷<��?E9�T��p�<���b�s���`���=6EScu�)�>4�M�O���F��j����_�<
�0����F�����qd&���T?C�A���Rˏ�Vt�Yp�s�kɓ[����pj��,AX3�> �bj0�!<���S���.Yʊ��$���M���6�{+jf�op�_Zq�g���\�-������o��u�|]�E(f�,��I��~Y�"��A~OQ�Ӥ�m<�=���̂�i��Wf�	=��!���}m�  ��6t%2�I7s�x '��@-�E�vQ=����Q��D�.�W���5��;� Ee�h�K@���3��Oj��uM2�OO_����uԈT�l�Ag�hX���IM������4���N;�.DP�8�I%��_0'� a�܎��TH9&��2s���,������:�\dNé7$���\��2-7���1@6v��q'�+�� �a�]+��}А�OhS�d�I@5@2���$W=�"�Y� �a���.d�^���Ǎu�a ���4%Sst쎓�MOST��$r�Ƿ��=6Q�u��ek��
���!���x=�o8�u����o ��(Hw�hDip�M=���@��y+�z~u��f�����J�9c��+h�"�9��Q�T���s8��<�>��>%L\;��S@k�JUS��"E�AO��:+(;��H�����#J���?˻W�Ir�e7�u45~I=�ۅ�J����HVo�#�2N��T���i̺6��"�U��T�R=�\Vޛ�U� ��	Rq)�Bm2fΛW��e��p��e�]�U���{ɖ0־�<fR���ntÍ�j��o�d��T�Ͼ̚���6���'�dm7�'XA�e�N��7�.f����a�,;m���0 ��y�r�D��>wL�䩒��a�R���-�oq��&L\��@���e����◌�Ɖ�7˄ۘ*gs���򜓥�R�Fޑ����*m0���	������nO���T)��S����3ak"?�O�[����A&^�B�x����𥳐��<ިx����h��z�HX/yi �W�n'0�&�n�+�r1O��ZrUk�&i�e*���u���u��vXF�PvA1G ��̱WX$��*d3_��"k8�|��w����P� r�X�V��=$b���Z�}�6J.��09^<�먩����`��X���˔ҩ2K���Ƌ��>��Q.�<�-�fz��=�J�Iu�"�I,S^mP��{x�a\E�J_���۲ $?Ĺ�?��߬3(��$Pβz�G��zS�V������[�'�_�MY}����_̵�U֎_Zӯ;��>w1�6��=��*�"�=�{���要 jcF�0C8�1#���.&6�pOc�%`�>Xn�H�6dn��?
�+��,�#��i�~Mj�$6�4!g?�2wd	G<���P��ր�8�	�T��I��m
 2����G�E߁�  � �f���,t`����6%�C�h��
�x��o��x5� D�B��2^#h"��������Rd�)u�	�6r*�Y7�U���Y�1�%�ҁA4,X"��s�L�M=IL.�/��_��