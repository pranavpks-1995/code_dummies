��X�)�6�����J�S�y�$���GI�ԫ2p��ӝl�q���@qp.�P,���GX��_��ϥ�G�*�ăqHXr���|�C��e<��Ep���������!��8���UXȊ�+`�X��T&��a��|�i��¹��\N91��J��f�ؾ��l;Tb.;�O6)	��PQ����VY��S��Qkt^��rl)Mu6�n�E�@�	u�~�z=�I�'���{]4�.�Q^Dw�4Lh��*���PIS�!6u� �>0[j�cE��7i
���V�N[p   p!��9(CUT V)��R� ��J��3��ec���x(����PS�쭵mXW��"{$6�wY�F��􏿇����*|(�k��@g��Ɩ92	s��v��(9t�:��kVrx�T����	�@xlA�Q�������NI.��Z�����oi�z���� �     p!�Db# *X�-�mx	��K#�k �ؼ���� �
�቉� �o-9d�����HYu@B;ٝ�1~6������=u_[���|�0C�ѫ��6����>�-Ju��6w�-4�(Q&*��V�D���n���0���m0�n*K�}���\w     !��F0���D��fkB�r��M��r�Z޻ł�W���3��#-O�wb�O�pC{�J�om�ka��}�����!|�����W}?��k=���\	&L0�D�k���/_�
k��A|~_LO������ ���]������ꮣ�_<�� `    p!������B0�\ԗ���i�_�� #� �M7��"���8��$����Q�OU��c�|�a[��!�b߸kˏ@�?�ן�xnz���m������k�{d�Ą�)N 4#��=N	>��Z�l� 2B`�0K�H@S�.s����� !����1�H�! �R� X/G��ƀ  �#A�o���{���pA����[m&�� �aV�Q�kM�`b�^��n)N�o�[���a�C���`�����ф� �f�p]����>(T	B{��
��̠��a�1�  ���z3��i�ga���e@  p!�������B�
�Y���
�������! �~�o���LK�9C��X� �G-�_;�V���0���N�#R�Y&.j$G��b�1�����";���@?�����D|�z����Br.H\3�P�ٓ|�ư�� |�H�;����^A�0   �!)��E�Ca�,��ܻ���i*�,͂rr]QdD���0���p'H(�ݓe2�=�V)�|k�����ӑ�
`�pެ����bJ��I�F�M|&�1ޓUƻ����T.��f�_v��MY_�i�?�q�{k
Gm�|^=uR����A ׳QL�D�"(�#�! ��+�f �I��˵ �j��`5i�M��A@  p�K��=   �Р����C����׭8x�ڄ���R���]�h) ���Q�A���l����z�)N̡p�'(r_+J�]�����`�\�}�g�3P�-%*��Yz�:4�p��x������m���q헅�3�6��5$�'+\nJ,ˉ,������}���=�R?�0���%iGJ��p�J�b�9�: e�x1j	�ڐᄀ�}��D	�=m�;*͐�-���n��ڑ�2m{�<G�ܐ�J5��H��;�����n"_k����h\82�Ä/�%n���D��5��ODtlv���z�%X���''��sy�{�\�N2��=��J�M��,���n�O�@�=�2�bι-2|1���[;*�h ��TW;�Pk��Z�mO����,.�.�k��HH����g�YY��'���M��4y��
�yP�o#����H]���g��`�(sT�e{�.=��T�0���[��k��^Y
�k;�����J��U�I�TK�v?���L�.�W��C����M�$��j��}�B�n<ȯT(陥�F���=�Q�<ug���6SnE �f�g��U_kko��Lk���Ҙ�'�	��}3�e��q�����B'�e�?�A��Iڙ��Љ=i��4�U�=J|�3i�"����׳*��@��v�i���+`�!�,<Qb�Ȉ�U�B`�:��)gs2�	3Xx�'K^�䦩�HJ�=�.FE?�~���L[����!��<���N�������3��O�ݝ)���)ۿ3�zN�k�^v�jt߭ޢ�.�~*Mq]��S7��\xܘ��*���e%�|R�m�� �r�������%��:������vF�N=ë�s2W*bɮP9 o�WFi�J�b���7�}�����y��[xz6������m����̫�a��j�	W��������X�J.��f�8��W������腒>�yc���>	���^ו^���]��T�n�����d���s8w���m3�P!ǖk���O~��$-@Z�}���u�qX�0I�S�d�|so�wT_�(�	��@+	`�|�{gh�1�E�,�E�	�C�O��@"�L�F�*_6�x���G2���9��3�F݆ic&=����#��D/�Tw��f�HW�ڟ��:�=3g�M�"6sV53)�?����U�β���?|�kV���o���2WЃO�4};[���g긪_�0��9�`�_Tѽ�7���,��y�֟�~à6���v�1.�&�W��q�@1f�ꉞ!�ID�cr�S���*;n^*��]p�ӣ���٩�
�MAÝ��S��� x7Z�*0�]�Ӥ//M����I�Cg���T7kkq1IW�����R�Y,�K1z�L�__w�e�jU��(��"��#���m�$��G�lZ�����`�32�:h
��߄
6@i�!�3��6 x;�.�tQq�nuiʳ%ڙ;��v��R�K�x�%�ȫ�r��i��5w�N�����r�4n�7ߧ��(E����	���;g����k�ٶ�"M!)(�`��>�3>�䯶L�+mJƱr�֐ȗ��0���	�x:�����k?�ͣrNs5�1{]C'�8ɖ�U�'2�}�i� ��@��G�$W���&��*��7�X�6��.��g���u�*�ĞA(��$�F-࠻�BP�ҥ��V��z�Syg��k�����_]�G����&�m���D�q�՟PB"���Jh����`���ɒNFo�=�S��f�B򋗾1��w��0�����)��z$����֕��n��f>9p��縡K�}���NS��AV%��ݤ��mt��KڋCڥ2�.����!J��q���#Й�9M�C�?H�P���C_		��?@ʮ%��<)I��Q�i#��_;��jb� ��m��~w�O&���s�����ާE0�6I������n̔ϮvB�3��_��