}32��e�z�m���S�
���bra[ʏ<���"=���x^���t��z��y+,�NG��]l�{_��8lt�8�Μ���`�,uP�6��9y;���1�u ,��V�6Ϋ�&ҕg�3������#����N'���9��*w�=IQ�Ur��cQ�pcF�[67�C#otA�pU��!������S2ĲJ�4}EĊ=��}7�4D�ހ��;;�����&�(_���Ϟ����}�@�h��_��4��C���ݠ��6'=D��#���Mľ�D��ሿ���L�i�B5$(޳�=�mq	7b�>��T1W�J&9�>��������b��.;ƛq
��n`���䵺y�����9�[�p������d4?�~���k�s�;0�]��=�uI�%0����
�c�#��D�� !UQ���G�~��i���J���n��|��eE��̔�H�I� {2P��ooFB�?�'D��Z{,�u���e�L�\�'��*I���~�2~��1xޢ��g��1O��J,���.�a9CB�d��=MZ4M�i����i$3��!ޯe`�Q��Eo�8&�l\lU�?�ɳ�drb�q�T�瘡; `�D!У=�z���͘��� e�����0�Fi
U!��Q�|��>K�G�u�S��^�(���R]�jxpS��'�A�i+���Z�=�U/ƽ�<��6���p��G����o�j���`i����e��Qj~�
�ѠQ�Q���9�1.��=�^F�C�(\��b%�o
��D:���i5���fߓ�� �A���y�'��@(��G)Z'��3�5N�Q�������z,|�D�a�����*�!i!;����˭����BlC
/�W�����j㠴��m�JQ��Y�������"G���Ud��S�s���Q�Өӽ����ya2n����H{A�)5d�!&��7xg�`;iGɡ�X���D>x兮���w1�D��?,��j����d�K5����^|ћ�������*=d� ����T�ܪa离՞t��௼�Bؕ[�H�$'��0����b�b��.XG��-n���sv$	�{)Y>)��x�e����x>�+�1en��yܔ�=ѐD	�<��y�c|��͞Q5�:A�/�����%�$`}Q�j�*d�~�n<��aٓ޽1����.L ��B�9��iݭ�*��K��x���+Z��9�ͳ�&��]��|T�4�ɲ�q��5��y�<jY�$�?9S�N��;ܜ�C�H�,��4Ⴝ�`�C~���@� ��UJ}���PǑ�n�:oU9�쨃d0�m�ڡ}&/�+Q�x��L�V�*Zd�r��/nW�VL�'�4/����¸a��[ד���B[���4)�̈́n��'פZb���u�Og��/�M*�wp� J@�m�N�HK�����MFaM%	�g�J�sh�N`�G��X�Ӱ���ң�4��H�JƐ��ᄰ.����� �f K�AE��s��1���/fFS1t�J�Kِby���5t]δ/�r�0B* tP�{{�������3g�ȳ�z�q�2r1�$��ʾ$
��}�0E�A��W	H4�F�r:V޶�L��\N����H�YʌT"����"���5�-� �x� ���ϊq'�u������H&��}�Y��{!x��/x��GNd�e�aw�p��Da�kҝ��~O��Fr��v�ho�������	�~X (��G�(I=�)�0��=�?X�m���\`22�W���'K[�����z��R�
~�s��a�{�I�+�I<ĸ��94@�	��I��kI�S�n%�I}�%��θ�Ϙk}P �9�E�=�