>�V�)��n��G<��������,�YĴ����Aܫ1�6�=��[�^���d�S��Az�Q��#Lû�ìӥk����S�n��݁>�j�v��'���֜%�>IE�t;��R\�[Q&�a$&�����yG�l�`�w�k���Sf�w���U,�Lͨ}7�<�md�ψ7��ٛpR�G"H`q���9�v=r�#��S�~+�O���GD�g�������!� ������?u/�!H'�d`�$��4�k,ھ@iء����#J�[�Z-L�ɶ�]���n�A�[U���5r�+(�	���E�B�:�P]�,�d4T�P����6��
͗���a�՞rm��|���� ����x�I�d�}A$va:7�5�ai�y��&�F4�$L�t�%��/�����LǭL��^�k���ԼgH�ȩ��ɯ=x\Ջ�Ķ��~bsZ0�'嬫��3n��Ru^�u��ɗ{��P ; ,=���y?53��2!�"�x��r^G"���p� �@�ڨ d����0�E|�F��hL�a��k͈c���D�
'�N�q�0�j�#Ut��i���m7*��1?��U*��zB6��Z̎ւ�w���Oq�xxR=ZԈY&[���Ep�6�f�w;g�4�](�� ��fX}�9�e��3��V;���$�W�[pAĚ�&���F�~�Ť+&��������u����ӊxw�|*5�I�=P5�3P62f���%��Q(t�N���pg+]�r���uo**���1J��=���˙�{������+ҁ�}��u.j��66��'��ޓ�ķ��кVTm�-�n�l�_�M�2��h9q�rъg�ٞ>B/%N��w��ip7�y��G���������V�Ҿ�!ñ����jϒ��b\�JJ�d[<�����D���V�.:��vGm�ϊ��9Y��<��kzю@���o׍XƩ��(��ʰB^��@
�е��sVXn��Le�����ء��١���#,U�lX+o��wE�=�ݺP�EZL4�ES�f���h�~�o�a��.������繹��&4��R��QB�%�ڍ�!k��7J�(We�s�M{��ϹOk���k�86��.��U9E�r��#���wm�B�	����z�gP�8�ඃ��z�U���j�:�Q@E�qz2�d�2�"����WR�� h=!A8�W$��j���}4�ȼ�����\q��N�p�s�\g�{,�S�d�û�:�"$\�[�>�����w���v؟+�����I�͹��z �	4C8�_��Tj�H��|LƜ����*De;j�5� !+ߘG��jm-�60�������C��#�3E%�>%xK��k��H���+;E�g�vv���β%
�@�϶�6ț.8����U��F�S�>���R�ۗ�=;(ИCf@�Z��*<�W:פ�M�A;��ξ�ci�CH(�ܔǳ��{]?��h@��h��������RK$�ƊJP�[��c�����$�oYz�a����@I
p��9�%���	-z�{����D/��MC�S�|
��B?#N�AL�	��p��<5�n�l�l�6���2@*l�I��q����㙭QRM���,4��	���g��VY�?�}���#L;��|q�P�fp��^Yd�3`t&��U%�����$���2S������C�dw#t��w�v�����.˃����4r�jQS*���o�C/}H��9}<H{/\.����<�fe(��J�RU��-x��<�ҍ�[��N@b�d�)�z]���C�VDasl�SA>]o�`.�_��m����k���+87��ܦj	��uD�K~{.����t��,�˕��D�����=*7fбZ�k>��j�jhH��i�����.ݡci{�� ƈs���Q�w�	��E?H�%AL�!aR��X���b_x���w���v��T!%:�\�b�T� ����H iRZ�V�X<Fp(�jtb���zA�����0B���/�{ g�&��M�Gj��ta��C�L%Ѭ��kRA���y�3�sS䱪i+-qq�{�i�Z;��ޥ�ZN�6�:I(*��ʒ��Os�f��V�"�m-��ĭ�'6cL���;��EQX�ڲwS�QS��*�h?d��+w�?ٝ�}W��(OH��:9����1�������,qc>���r�:h�Wc/�4��y~8w����װ�E��R����l��ؗЙ���P{���\U4�BR��)Uׂ�B�'p��|!�,��ɀ�p2tAp`���-�!�}��\F�#t�{HW�P�{��$��+��a2�h�QK�#���ئw%� �iBy�$/��a�H�f.��t�ԲuVw'���%�D�f�1���cȓ�?'�.��oD�����>?��X!����]ȳ|V��)��J����*���e�q�SY{�yE��%�����ͤnM\C��O�ՈO��+Ky�n��Nx_[{��	0b��� �	6��Y!�������ԏK.|�������
���6?X��y�d�R>��٧�_��a
������W�;�[�0�Ȑ�����;n��BxDG���7����>�g]�`A�s���Č#�"$����{tb\� Bb��~7}0�����1D�Z��,Dˮ��y�l�@�໇Q��8�g��O�, �/k�a�8�gԆ]�5L@K0�%]��O��k
�|�y"����Gp�W��o�%�h���2�/3�8'�[.��$r���W���i�>��O�":L���6�.�,�#r����{e����;���`�~�S�͹��uŦ��z�����x��~���*�@�rK��Pڴ��iWTc��b��X�|{�g�8�f`�F�㣞B�-z��\��b)&〪��uAS��Q5�È¥�~�� ��� ��iʀm��6)�K��8e�-�*`�[��@�f���"A�j��ˋ��;�r.4��Y�n, �j��}1%����f�y����0"�]L]�ՎZ%��ˡ����O`I:޷vI�r�c\��nGe��}z���R�UI�Q �a8�z9A�Z��r�lH�� ����9��!'m�>��l>�E&�H��1�����a�����p� �]�8�P%y<n�+e�ɭ��P0��	R܇6��@���}�3$�֎�q � A;O�_��iV���8r���@��
_$;hq1F")eݺ�!�.Z��s���Y��I+�ؼ�/ ���6�ưGEϬ�*��mԪ �=d�Կ��C�q��K5/��i>�̵/�q��*?�e�F:�qc�zw��46%�h���rLk���x�f��E��s"�۲�h��f	�.Z0�ATC���'��S߿�zޥ���{�[�onǂI1&d�X/J��u+�I�Pw��������?z-��T�����4H�
�-(�npw�i��Ħg(�W'���[�2~K,�X�Pd"���\�J'�j^�
$$}+)|hY�fy+]��zs��#�p����%��f dC��,?>�0熐�eT���r��ԱA �4��h������V�?Bҵ���Б��e*/h�Y���]6��Y��f!8B콿z/7v `���h�:h7���U�!]�����@�g��m�T1����0��T�nuJu�[8��f�=�"��W3
��w�	�R�2r�\��/�����cι���P{�sp�D�i�SBK�����.�D�KՒ�ӆ�Y�"n&���tG
<(�b��k߰��4�Lw��S���R��;�)�;�����?�_��-��aXY�Y!����ZO�����PE`�c5����x�@OX����@D�&�G�Þկ�����ϗ]E'�L��k5a٭��Bpf�W�} v�F��'垰;.�&�d�u�$���� zB4xVSK�o�M0�Z���Y;PrtDj�� GT�{G��p�6s�Yͮ^ց¡H��.�"dE�[OD������E��,����ZJp�>T���tͅ��&�w����B����o��pr����|��(�w(b���M�)�;k�������$pv�!�*�d ��KC<r��ת_�ù@�B���}<�9��X>��j,�v�g��ZRH;��Y�D�c����i˷�հ�Ӳ�G?�}s�W� ��*�_�9"��T����b�1P�t�*��fr �Xð�H��a�;�m��P����̀-�����)J�$K�1�5"����J���C]�*MXee��zυK�U��?�O���o��KSZ�T��-�bܷ@7�̴�-S|�ΌW�A#�xY��T�({A*-+F��f��]�FW���\� ��;]�C�TR��J����H�SGpW����KR��Ȉp���\1�aɆř�2έ�ָ2!+RG0P���c2oI:@�]Ԕ�ߴ�����)�2Qg�����I��=*R~�1�9��]ά��	p�A�
������T��eO��.�QΒ��HU���v�Ps�:�w=H�����_񥂓s9�A%�]��/�0����w��q��.��|}늓?�,�^������צCm����� ��K6��F�� ȕ����-*2快�.����M*ؙ��C�n���N��͞�����={]ZMϤD˘��Q�����4��C~�orQ��ܼ��?"�q�����S$�O��I�'W�C��V['r`��9�$&�?�"�q�V+7��ͭ��de��f��q����
�n��R���ڿ�Eeb^,A�}�} 6&�d]s�̓R����q�g��7õǯOn?�%S�x��8T���K ��b�P&�}{�dA�#QE؈� 	^�/�Jt�����~�'�rĀf�$��)��s�,��M��]1��(�L��P����X�&����XjS]a�0"�Ԕ�޳��b��,;�L�l��;lΙ8���b�hapM�Z��<n�%CmZ؟�1�.t�k0�;ds'�)�h 6�������^A��o_�	���0ц��B���"�*0����x���tb���c����8�	�t�k��n����Z�ɉ�=Z�(���b����lGƒ!V:�w����Ǚ ��&2/��0/�t?:��[ ��?d��ޢUڷ���0����很O��G�cb���5ȍ	!2���N��F���;�$[�?���0.:���u���A��3��˧Ȝ%��g"����}�C����8\M�V{�P��}Uu1�D�;������f0�~�1q{�j+TE8[sQ�c��u}m�D� �D�'�%����i������aH7���)� R<�G�������*���낋�)�B��x��G��:���,]Ǹm��Z��WTϤ��}Zʡq\������VX�uGaN�ْ��/8{��[,>z
�<��U�q�ū��oH1��|����+B�W*'�h��Rm`��XGc�-.xN��X�~����$�C�����D (N��I���S��S�q��+˴�N��+M�hV���zx5��s`�䅩)���pyv�Z�S9v�s�����	����Z�'7LCj��{З�J"m�4&,.v�����Dl��G�E[��q�0+"T�N��� ܐ�[S�$p71�?o�����4	Xۜ����]k��,$