import BRAM::*;

typedef 4 Numchannels;

typedef Bit#(32) Addr;
typedef Bit#(32) Data;

