����;�Vr�L#Id�T�卩`>5?�P���1��C�N��a�^BK�/u�H��]�D�D��j�R硦��K�������R��WV(����n�'n�-�~�o�\cF��L#�N   ��W��c�F�ި2�H�!	��+�3��!�	��{o�����w/Cז���\F��+q��t��t'��t��u>;׀s�fC�.�i�"9�և2��=�瑫��y��t�w�՜|�o�7�r/t�f̩���0;�,<�3��Y����F�e0�30�Z�(Vc冂�_SJ!��~��5��,�<=�Q�L�3��i�G�۸|�nG���1n�*�	�js�����~/������S�=�#�.��C����j�-z�69�H���.���MJ�u��/���!����k�jOQ��]��2OC�մi/�����,ܥ7��׉���dTQ^�i`���C����CǋDį��+�EHz��uߙ�K��w>��B2����t䷌�Q��Ao/�<���J�N���"F�$��An+���t��sx�y*w^;��QR�;?������Lb#��F��f��,�g^Q[�� ��kn�6�u����@n�#���r��J�>��9��D�͂�Bu!ƚ�'ѕ]K�t��r�8z��;߹e�����)v,V/��w;ei���y;3�������D"� 0��6�e#s��s{:��X��?����z��� �#����.��&������:i��Z����`Q��Ŗ���K�M=�B+��c�Ͱ���-����p��f�u�ңWY��/
��PN��O%O����JU3D3h��&�Ο}�4�o==W���v�o�w���;��ɞ����)8Fi�{���,'�H3/U��+X���0��#)����q������Z�0Y"�@�\!�4��Wx���;"})Z]�MP�S�wD�49>4��i����΂������l;21��j�1�PH������aK:���U͈5`�$�.]��x[��������kZi�*O%�!�P�X4��<Y�2e�����b��*ƙS��׵�{�͝v+��IbP}���@�"v�{��y���[T�������幇ƁF�|p1e��K��ǵ�3��j��N�W��������^[r������H�ER�es�=�\�<�hU��Qz��O��z\�5�V�NZt"70p�7�ې�)���
h��T�H}�ǹ7��3hh,s�0ͤ+U76��� x7%0����~{�O��6�" 3�.#�u8��.�b�w�����̨��1F�;��e�!�k��%��i5A*�l���0(n0����a�^}O����JX��������d�!������}�7�����+���/�!�ر�~����o]c���Ɠ�r��z!X�*�S�%��o,*͖�$�]��������6]o8�ؙ&t6I��ؔ��l���42��;>�x�6�F�3<��˫��of���x^�%�u:�dbu�n����%o$�k̮�,i�d��=��P;u����t�t�P�7�{B�ΈrARQxK�i�f��V���JDi��Dd��&�{����wF��*�:[չ!�����O��_[:0��M�J]'� ݂w�}�?������<�S���W�$���NQ��^�O.�����
�������μ)�o#;��4x�7���0���Pf��k]����(�FK�bcSu�ҳ��*a�^B���C/���-���W�����1|r(�K$����ӯ�D�ʮ_��H��Gk�f
�o�yhܯծ(k��{oi���F	W=��X:��d|�2������if��L���Ǭ�(�V��ҡga��ǩy�`����v�	CBי$�cY��f7��G����F�=N���̅��j�4(Rj[��j��㦫�ƣ�#.p�E�E�l$�8�56��3>B.������q�O�x=Ʋ(l,����Q��G�n�ӏ�����'O"�g�l�)`f�����Q�mY;hԞ�e݈Q\���0�܈}�(7T���xuavo�H�T��;'2H��3�$����yC"���Z��3�U�aRl{ygj>��j�8P�v>�/���8�3)[}���L�����F�̳�U+O�2��C�N"���GD����+/>�M��$���L�Nad۪)�ͫ�H����^����K�v[$��Z;��D'��w��+kL��}"F��V�P��uLf��ߧ�R]���� ^:"�e�bN�M��/��~6S>7�{��E,1�Τ3�O�K�E���I&oE��l�������_i��n�X��[8���ֈ��̤�X���f�d���#���K���PZ�̻R�4Qm�͝�h���踲�g��r�(�45 �9ԵF���mA5�5'����v4����)�x��@�a��m{2�ǙM	��Б5W<up��b�m�56��R�9���ط��2t˖�R�bX,�]S�*���3���W��#��r��:l^��h�1�z�ū��E+a���Ƈm�@�LB�.�mO�K�Q����v��/j�m�0#���az�U�����m�d,h�`'��q$�Y��b=oԨd� �<71��Q0�'���vn���,���������e��|��EV�q�p�������^���aP����.B=�M����l+�m�q���۰��R��h��p�'EЮ�� =�0̀��C ���Ce����sun���2�v4�������.=p¾��0�,R*��\�s"�#�؆zt�l���-���9�*�a|������'�h�)��*VХ�Y�S#[�u����UF���
~Ϸ�8�oK�N���E�}J��:ۙo_�F>SZ���K�n��7����������4�wd���gPle �{��dL<I@�FzT�J|����rb��H��<T��+�K?�}1	*S�MY~��˭�ώ�G)�cX�`�T~��W+ەG�*tH4�y7�x���H�ץ�Su�>�\"
�Rh�O[P����aK�j.ەF0�5y�>R:��G:�N�0
=�*]��tz�Uů����E�[;�>
5������G�s��t����#b���]�x�mi@��`JL���fr��ITܾ�?�@^N*�S�X��4���z8�b9֗?1n�`��І��sI�o���C.�$  &�"%W��:0E,#;� ���Y������� {_����Q]PO�;��4�}�H?����n��U��������FAqL}U�'B��9�O��BoAl�ڷ�9pg7���x�q�U0�	��`�<�\���T{�_��-{y�&oNg��ͣԝ���15E�ń4NQR�B�nn@��<�@I��D[8ۿ5�l�JG֕�jYM��*Y�:��U	���=vdBEs
�3y��1� 5�����|��o�>'S;�#f�2Uv�*���QQ�hPN𳌝��ȖH��>��{���g�$ьp<����Y��د̄R[�|Z1�V|���W�?��(rQVS��Ά�m:��;�u���u%D3@�y��h��5QKv$$��/����`c������w{sV5�_�@�n�'v�:KJɀ	z+Vگ%�Y�٪���}/�fdx'��,)�N�5�F!D2���N�o&d�=�ՔV��G'}��f�84�dva��x:O8n늜<U��{
�ܯ}w#h�ښ��I�έf�J��U���b0�=Z����O-A!�\̈��H�3E1����ׁ��o��{���?�u`]r@�]ie8�QP�&_���@�%*����Zku����9��g�5�@HpK�tsW ��I$�y�N�	!���p"���?K��h�خ�{I�Ogh�!�J2F�cު��9��(��oW���9�H�p��z��Y�
;�:!'�6W;�Iet���f[�3���G����B�;b����56�����%�����p�u{��T-أA�� �  x ���H�ч��z�� |��$z����Myg�a6�|;3�|�7g���I��}�}�w�P����N:�Wd�>�P?4�1�R2/8#̗�ߠlYK{1;��^�.$EL�!G�F�g%�h����53d� h�L*�j�b�=ĭY`��i�ɏ�F�X����Rb�k]��z�AC>�����Of��U�΀���Y�-��SE��^�4ѥ�<�O����@7Q2�b��(��jz\g��:�r�q}
`b��t��f�C1h���sw���m�Q%�P	�b,�C�e$��h�`v�O��/� k[�/���@�X�P�}~|a�58aW�����I��JO�U&*��B�73Q��Gƀ�ES�g��������!�)�ʡ1HL1 �U�^t���
��C� "����
���]]|�_Z��1� ��F�.�sb2
���n���EUd���+���[o�[P.�!��P bڤ�τ�c����0HW�y��4Q���|]�Q�	P0Ke b�H0� rA��tڙ���$���B9��    8!���"��,,"KRh��V8 }�a}�8�F�:���8�C���9���sH��_���f�s~ψm���p���x�B�DZD�,��+Qܷ�*,�"���(��,��M��Fe(���#3[E�ɼQ��d�:��-Jl ��v�*�q)�
�0  p!����3�T`L�2�Z���W��B��D��-%�꽷3��/�~CB���|f��s�Pz�@4��<&y�9���TZ3֌�- F��w�o����h�q������-*8��u��x�?��u�>= cr�� ]+dY� ���ݤ/����9��   �!�
��ꢸ�HQD(
R�bXR����� �q8qj��&s��@�Nx��ʕy��rг�Sш�xӇ��,4Y�V�����wOgB��<�$3P����E�+��L����id�z读�2�<anۧP��� IA��B ��F�(x����/����(0  !��DJ�D +%�K]\�k~'�yV��(QfG��?=��?�=�{}v�a�+�'�v� �����&�:�U����ڪ�"��Meeu��9RFy��ݙ��&��.��Q�i]��?��!��ʣ(i@,�(A�p� $WB5WH�`'��X;�<ʶ>��!xM�G;�|�p   !��!`(���  9�%@ �NR�n�����;�I\���]�� M��1�����XJ�-u6���Z}6��X�t��*2�V��D	�xz2g��Y��Q��2��j��O�KU'�d�T֨5��XT��!�M�@L@ ?�� K�� #�+����Y��w\�    !��&K2�Xh!P� ��B��BR��_t��I �J�ҝ�y"��|s�����$B�����E���PJ�r|�K��-���4�������m��1�8OM:��H�")���wUF�r���}!k�0�0�[RHx���S�K�ʱ}u�5K10s�X�      !��
iE� �@� �,�a�>�nDJ��L��<�n��I�N~���s�p6��6��Y��K*Ԍ�dƦ /� C�by!��x��N���>���0R|V�Q=%룴5�MdY5�<�ONgge��w���\� �� S� �L1���n��듊)� `    �K��   ��0�u_q:0O����k�f"��z���6Sح�Μ8���E�0=��M�����ր^Z�6��._ͩ8�������x��8�V���S_ΐ^����
�����:Qj�4��S��
;oB+� c�'*���]�kVP��.�0?��vmzS�t��6]s�o6�ȇ`c0�z�D��M�߼Gm��wG|�w��`�(/�yж�rTF����_f���D�����^����z4���]�\h�7��~�G��C��P�A�_�=d��P�j��؅�	,�q![�( 01�#�tP���~��m8i�l�R�E54HǑ/�c#~D�}�]���t�|G��ؾ�h%�#C.��6�NǢq�*��:
��׵Z��&0 �sY/���G����;H*�p���10	�����Y� &Zߤ&<2��Y͈<w{p��X��0 H�yxLN�{��4����ߐI�_�ƫ����	P��_�j��q�ԫsqC$�Q�߄n� ߝ�:k�ŊP��UW=�7~��c�����Ԍ�'�h�Y�[DZ�#)��R-je�4���s�F������WO�9L�<�f����gY�|�\J�i�z�4W��
+�s\�v��8��u�n������Qn����=��o6r�/�_�>�q>��m&F`n1�  �{/����V�u��7���X[�ޜ-�x�A�g�����2ꏀ�Ѣ���e����n^~^9<��k��N�A޻P�+!��G��{:�)G���.��Wa���xa���F-�Q�hFF4.�sXv���*��������eF�����Qª��*��<N����%�oϠ�� �Oo+;j?�(Z�Y%�R�|X�E�ir,�x�ꀀ�.[���]����}|�p7�Y,D&[CsD/����O���ү�Wg>>dm���]�^�Q�W��� ��{��L|���Z��Sb�E�6w���
�i��" Z� ��G\9� ����,�5��,S���U|I�������w�S�cXL�II]P�@�:��e�*-~v��yyΉD.Rx
U��@��WPT��t	(�*�(C�.l8x�%��݀#D���e��v�|
�����V�J��_a���#�/t6B��>�ES�3v�;S��i\ע����}�;����_P���Y;'f�6ˊ�w��5��+l��}!3|���QH�}�q��$.�Z9�����`Q ����&G��s��<�/�s�o��ٝ#�	�]�g�E)�{�� k=����Z��BG@0��q����`�.��k���q��>c�F�с���D)�ѥ
seqCb=�g��UF�c��N�[|�j#n���H�L}�T���bJ-���9��,���E|�<�w�!/���J��#�y.�E$p~�zV����0�W�P��u�E����[WK-o�w�����l留��Ґz�.㚅X�߆a�𢬟�>��e8�|������l�b�'Rߩ��%�A,Ni~|F���B�e�����(��'���y�!�Ѧ��T�F*Zj�&��}��z����F�,�F�^�S��~���Õ�K�`j/d�3]��� =R���N�Y�q��8%?�i�`�(�	�|D�=��Ac�J�i����Ѷ&�{��1�d��Ļ�i�*�����R��7B���]ɼ�.)�7TKW�l#7BKZ*�}�E���=�N�Rtg~�!����K�P��%�(ݗÝ�y9b�P�n��^�7��V��q���s���v
I:�q�є���>�d��G�A��q�RD�� ��K!͹��ᘓ����<�r�)�+I�XM�%D�5e��S���M���+`�]�G�u����yр��s�g��!�ŬzT� c� �{.`�F&�k�-7��&�ZL>��f+n��T����g{�g"Nn��D��s��3�_���&/	z�g���ˁ�"��^�^Ex���^�{���Fa�q<�S~#K��{[�4%S-����L'�r="��	�������J�юU_�N��N�M�3Z�y�ʢ�6�
�zʥt���TF^�{�"��xq�[�>緰��pC45��n�Ӈ29�'�o��f������& ��;���@=��`�]N���vB���ꍯ4z�6�M`�4x"
��&�D��/��ZU�DN�?�I��N��+�Z����`7�]u���uK���Į�E��*�,/F�a8���q�RN$p�^&��]@�?X��~WrwQwۺz"�׮ـ�y���D �
�H
��2��(V�����b�&��Sie�����J�KeF���)j��7B<�\KglG��ՔNr%�Ni��[��[�ta��q�NP�.`_��t��b�0'�a"LOF��Td��p�q��NQ�Bn?��E{���A�`�#?ԧ�Lew[����5��L�VycM�I��gF������`v>ǲ�F�ָ�I%��_��c���fWUfi��q�/�R3�@��%dӗ��'�GkI�-��gw���^C������g�5��0��0PƠ˰�ռ,t�� u#���snH&TwF���AN�Imv��[�G�3��!�4Z�0&~���6���̍x������� RCɷ��;��,K��T&c���zԭ��A�(���t�|z��d=�ipS(���?S(B퀆�b�B͢a����-���)A�����b	���*�b��[��Yz!ګH��?y.H���Fʛx�����pH�EXe�� ��t�i��bkxF��D:�r�\�OjȅtX)��/�eԹ�y��J9[Vx�F�I��X+IѽQ���]�����T��@�uC��f�	��&3�E�y���P=niD�}��N��_ҫ�v�,#�;t홵���	�����?ʍ-�� ֭uԏ�k�*�G�@˴ws���v�H�BX%yz�G��ݜ��M=X$cB�� Q[����S W-����;ĕ�#6����E��7��ѕ�'b/E�T�!�ޏ�����6�\P�:��*��� g� >�*�CN��  F��%�_q��z�ֹFT2$.7�6�7堧����t�h۲{F�AA��N{��/�쯜N4S nT"�=s�oĴ�(993���B-1���7��DP�K�:�b�Ҽ\b��Y�6J&6���a�A�Et�?d����ס'�TP������t�)�@��o��`l�پc@���W���Z(�V�M%�Fgz`�d�<���4|�M��T��V������@�w�v?�F'iُ�S6,�X���{�H`wCQ~ݟ�ƕP��-`F�U	��ߊc58��l��Y�@C�������¢�z��@��^�c��#!���Sg��|m�)���w�'�*=�l�ȑ5Mˀ���	!T>���T�����q�%C*��|��n��l1�c��"�!ͭ�$[��	66���\��QC7��4:��l�!�԰D�G�}���dX>������wY��%wF��v�&-�VV��f4fy,l�{��z��?H?{�
!4�^�P.j}�P�2���"��[:Y{��I��+��O�>��h�I�8�JyvҠ�i��='~3TK:�EwI�i�K<��J٦-U87yA���x>V�s�,4��f�Ti��}��Q��K������'����[Y:��Z�%I�_(4!�ZI'0I��U�ǍU��=R�<�� �KF�b��LK���6�2�ΦٓL�
2t�Έ�2���T��I��w͚���
�A3M��<[G��G�.���
mlT�)�jԈ������C�d9U�3hYA��պ�@lI
�`�*��@R������w�>���j ��՘GF� ��}��7��K�Q�����A}�x  u �f�_H�ч��a��0���o������N�ǖ�F�@��輢L��A��bF����?N��B}(�'w�Ck~r(�/��u����K��_������oj�1���|�U�"/�T=q�n��4y�,3H�RM4������.�SI�@��/I�i�:�E�����k���h�� Z������G�y~85�Z*��sd�_�w��$�(ݠ!U��(s�RV���:x���v>�kc�bi�.i�H�베|�F���.~5��x�
8�� 3�t��	�nx�+RT����C�P�C/����_Z�Ws?��03�݆~Y3�-Mw�e-���`��f,�EW��v���*��~�()����N	O�"��[xR9��B���Ao��   g �-�c�I�r	� ,H����wɡ@F���XY?�w�j�~>�E�b���v��w�~�w��������Vcw�S�s�6ۜ3�=&E@�D�c��a؇}Է��\�]І`:��*xzrT��g]����1�-B�<Z��}���ƕb����b��#�ȴ�I�3������b+a�8.\�/��F�ri�Mr#�ϸ��:I�	ֈ7s�ⵕ�,��`�5on�^q�fe�_��T�9.#�8g��9�nߴ�&��$*Ut 1�+���W��Ň��u�J#r��ԚR������ņ>�m��W�Ŵ���l�e�a���C�]���se�Ý̦c��`�J���   
��P�Uq:0Nۋ��N #	�|e�����ۆ �&_���C�0ۍ� ��$^���BU?+��ʠf0$��r�Mqe��/6ǟ�J�̱�blB���}�=�́jbB���ǔ�h��u,�'�I�nf��}��@�K����s3�_����G>��4 r C����{Ќϐ�-���j�-�������;V����
�)��b���^��>_f)��?g͟#2ݬ���"dp�2O!tJ`�{Q7\7�7�" mQ�
���~�a`��V(���ߙ-��f��R��D�U�f&p8�VG � �B����SQ I�X[F�ͣt ,+�� ��*t����d��H��$-Z����\;9>�˭�({�ä�m�u�Ɏ�s�s��ɗU�����R�����Ҕ�.��U��rDG�;��L:�N��9��Y�tH�C��Z�Ky�Q8�ה��������G>Q��j�#lD�3���G�].tA�Ao�J��Pk���i�o�y!I�04�Xh��T/