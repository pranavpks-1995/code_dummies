X�1���?}t�l�[��G�����[]�=:�ʃ7^Jr@�g �j󞷐��������0@���OQ�Ϯ9!��"�]Mٽ�!E�H���   xш����C��8�;�r�I �G-��V]��]��h�d�*����t��PQ\%��7�йE�AD!x�_�A8�s����XZ��8+���6���wy��dZ'�JKVs�]p^�,be��
���R'p��rzŬlrg<<��VN3[�����Js�Ӈ<�`hG�-�}�H$�i��Ó��+,�*���14w1��Í^1~{�Y�~ok[��N�A�w��>9��}�������-=��C��U��.�����	��R%�":����f8�M+m�w�Zz=]�xR���P��t�/�mP�>���S5ѝL_&�N٫����=.��}q���{nIQ���K�$B �`�����>Z^n.9o^"�iҢ�E� `�	�-k�����,r�1z��uI$kk�+ �-���<0�1I\"D�|+E���C,��x ��;J� �������or�#�\��@ʗ��n�,�!���ޮ��H�_G��9�,x�[�	�d�&[Q,�x���ChC0[P�ރ/��斀�i��|�����r�/VM�nI9m�������f*W��z��xT�1ʌP�K��Z�.S������w��%a[S<K�I" �[���n���N��t E��)��L����X�	Y�E�R��ς�d
P ����|'-���cʫ������	��xS�8�c؋�g���o�NFa�������o�|�2��Jp������T�^7�u��T��eq��nA���B��&o��C��uv�	{�2m-�G<0\���g��r�eo��ppr���ǜ�=������]�疋�t���}�z�������A�o��T;��q���=�SR���3�ʏ�W����Vy�FC���tY^�HX����W��;~��s� `lHǃ�'�"�<7�y��k���u�����[�k�2��T ����Z��Zk|pl	�&dos�]/*��
	�i~t�A5J�7��5Xʻ�0�诋�d��=6�		��D�31�.��#��s��&˗�N⽖��k�|�B_���&�7m*�L�0[f�)�c���˟v��zl�au�=�{3�g�l������y`���?����L�bH���&E���* �\P[G� N�A�|?q�����-�L>\4�+kL�֑�g*�iu��i�Z<~n���#�F̓d���OuiU.g1�Zެcx�
�
`[ �h�D�[2;���A$<���({LWn��Dȝ��<�����;��>3oiR����P��U�ȇ�� �-Jv�~�M�X��b�!�0��j���i�
͹��Q	}��o�%cC��z�T�N+��׎G�k�!�	�|?3ć#�*���م_.q��3�~a@r�H�
{]#H�j|�֢�p�+�׫u�{a-7U�]��Y�N�ɵ�k�Q�8)N%�����H�M4J&�˙G�\���(.wQ�3R�Rfl�#� RU�E ��x��ܺ��k�&
�:Q��HpF �Lu�n����&R稌6�t,����ʭ��R�����kn�!%f]�S���O�r�}�\��\��έ�\�6����A`��������[5[	G�@�3��=a'���;QVwu6s�I1r6��GK�fG����E��Eai���bqh��}�k���i�(4#|���^]�M�Q�������U�,���5Y~	� ߣ�H68xE��z=����� <vY���y1��%9�!�X��1�1�[O!�@�Ps��=fpC�6���jAM���9��}�	�_(�5�7�5�?B���Z=����,��f`�{��NI�`BT vu��4Rb��O!������J�(��z v4�od{�ց��v��Z�B�V�x@��j�!��a]��v�j.���- ��V�|�+�!o�~�7��G~�U�9s�d_�9`�(��P��"J��L�0���T�\��d��ב�����z!�������}��ǛTiE9>����AU�`�r��I��L�
�(��4+��3���j��V�r;]�q)8w��4��A��m��1b�0������\$v��9��Oa�,�RM,�w�K�=]���7�K�6��/��@)�X�{cw֤������d�����N�-.��¾nX�����$��{W��Aف�  ���'R��c�MzEx�$ix���%&R�^�v�↭Uxfu��'��4�eB+�&h�r���y�f�����G i��d��Vt����ʠ��@p/�R�J��§.��Wb�iJHN �:��3LZ6A�؂8Q#�E���	|x��=�X&6
� >!x���͉[���}�@�/�������s7]R��z����,✥��:='I�Js^g`�G�	z���,q�Z��D����~�TB��dOӇ�,`u�!��<e�h}�r(����.������2?q
r�[���S4��`h��Y����4�r�b3;uH�yT�~A��U��0�lJ��[<Iϔ�p(2K+���3�e�9�l�6C<35�Ǥ��I�������A1�����<���0�
�Tu� s�L����՛b��_��ғ�Q-�D_^PI?}���	�3P�Ļ�ش��5@�A$�P   ��U�m�9,�,��.�2U��Ă"��i�Z$/	7 j(9���"��t���?�@�s�0���'�����cr/�"�]e.�݀&��$f�St����`�̇�x;ם��aȎn�=��!�Q�����>� ��Z���R�ocC�-�N�ȰD�AG&f�A��7�)&a��_2�v�]g�$����	�<A�mo�9�5�8V��9;Ȯ.��+,�f"�c��4ö.��J��VV+���耇��(D�e+Q�iI'bP9��PD�>��>�t`��(K����AD�y   < ���u�m,a�T,�L"��Hs��A�-iC�D��n�"��-��Q�����2�����i ޟ����0�ΰ��,f�R��f��sU��ɒ<��aɺj�s�3o��nxĀ����3<$8y�w��j+�z��0�F|���i��8�L����M&�%���6����Cö&������G�7�b��y�{��M�o��0h���ϱ) vq$����M����S8>oݘq�H���4Ɠ�_'~�/�x
=g����ֺ\kO?���'��@��#c铬lVt�V�nz5Ѕ8�:��NN�Q9��A��    � �-����d�HF�E�Q���g���\bq=dK�k��v���8��55����wN�)xRj-c#�ą%���Y
2��L�6�� �B�k� �q �*;�]'�� v��e	�� 0{�l�������l7��
y%�Nt�/�eK����z��B��=��$M���O�fJa�JǮ�_ʵDȀkpBSK�,�$]'�PlL0�d��4:���1󦫲>�C�O<�@cs����}��Y1����&p�En�	g����ĩ��!��	T��T2�訦ZX:��B!�!;�GE�b�A�(�p?�k�b��Zq����c'����x��/��U:C7񐩂#��Q��4���lSnp��fў�v6
	�s������ %����5�{9M�4uo	��U�k뻻��J���      �!�
��
b��P$� V �՚�ވ ��r��^���-�'9<	R���
�\��T�G��$�N"2���Ak]
�S`����v��4��_�*�����P#�xI�յ1�X�e8*=���`.|<�H�DׯM�.��R �5��:"�kz ��˓��!L=��2�6ۀ !��V��0�bV�9K�e�K��CS1�gꤠ	g2i3�԰B�H������?�c��2�5�.�������,P݋.�S�z�ł:!
���	&���
;�Lfq����&��Ժ�6�h��aˏ�+/��J{�|�yf��ғ<C�V9�^�!UL�N�9�C�`  !)���a�"1�uZ8���2*5������U�(*>�&�� �x�=М��NV�$G8�l����O׳��V��?|�@��Y�J���^��yF�_9�0��8}�
e��2H��ʕӷzYP���Q\�,_}-��	V!!�� A0�&L�, ޷�t���>� o��$���-�;� B
�H�P@`�0!K�L1F��I�Ma
�P,3 @�Z�k .��'_CW�s����זe�$k/H�l�}�:(u�O�C�|�.�|��&�{�P���~-��J�֘�"|0Lk��+-�+dq�D,d�F#�4�y=��=W�֑u�TJ+��DJ9-'�.��<�!UL!���@n�2�!y���B���@!s����9�����%p�љ�����D!:��P���֍�o�9~���+m0��o�4W-u����&P��h.V%���#��h�M(�8P��4́��/�~����bBг���VS��	�|�ī�;K�I5�NvNj�w���l6Z���     !���İ�1 ! (� ��{������G��)�/�5{�eZ��N*�^ilRK��!U�	a�˃�e6φ��f�Ye``�D��3
{����9 D���)���.��'��ݽz�V���R (0H�2>3����l~꒕5��T� 0     �!����6!HQ �.��K�O  @jp�Q|o�8�Z�!��ޥT�[�BT�t�1����/��%{h�oߝ�r_rJ��)Zu�߭ˆ3-�Kt1�+"鑂��Hę�g�l,#A+O����X��>�&���Xl1��  q/D�UYM#v���x���'� 0 �F́	�   �Ѩ�U��C�����U0�l<��K yL���*��ӥ���RǊ�N}rB��5�1�6S�����;c�89s$��
���.U�ƴA��h�	}w$t�i�_G왬�� ˫�hG�`�z���  ���/w�prԉ��	�6J�<���eN�,&�ґ���5{�a�N�j@o�'S�mٓD����cZ:�\-
��s� �R�O1|]I��?m��:����5�c�U[�5i�����W�1���U���s��'����nb!�sA��"}�OβΉ<�AT��(�]�)���< (��cf�Z^-%K���h�s�Ū��%�I�x���ϋ�kpd�z�O<i	��1�kz܂E�OJ��Y^����	�b���,P��/�9<DZ�Tj��Ǻ���xi|,�1��Y�V��޴��s�1s�n�g_���,���s�u��Q�Ȇݷ�y��|��@X����_J�o
���m�j�����38��[��&E���G#�7�J�)5R��,�lrC�%�~�KéM��L��;�[��úq�\����$�c�t�-�^�:�/��`���^z0��203ٕOfab���K���.��>-r��L�?q���HG4��{z�7��&<�dA��{�3�$����W��a(~jU�d����l@��}=ep�ȓ�d��� �2S6���г�<��}���p�������9K[��$�<��VuQ�m�O{�����u���\S��G�lR�����`��\�T!��,+(�),6V+M2=�f+y�IP�Eml@�������{i\^�MR�ms��ۓ뉩B����L��C��}F����H�����d5)�X�[�����Z''�v���cq��G��{�b�&^���f� �s�6/��Z 2�����cZ��K��|��zh\�����{�i�Div��V51hM�Ҽ��Ɣ����eŀ���d�c���6�J	N!�(0� Q��*=��~�Y �3Ɋ��=�@�بc"ʺx@&b'�:��(fV�oG~Q�̟���|!��1���86�<�vz/�mlv��[qr�Q���P��]��p�cWx��JhP��y�1��K��@!��]��t5�z�י(�Y�� Q[tI����l�3�)�������&b�L��(����w��ݨ3XM��So
,.�`�	>&��{e��OA%���[��]�B��B��u>�R���"�Ե{���a��i����x�﫱#*��/jt��n�lN�����2�n^\%�!SP 鷎c��"����dpzy�B/el�>Et���d,f��z�*�䠳I�+��4 ��Ob�l�,4{{�Տ�Ԣ0��:�0B�k�_]6��B��ЫS��Juv���의����B|`=ʍ��x����?
V��	:M�t��L�b8��
j;NqK�5� "���s�h!Ng������O�Dwךgz;(̼�N���Rm�����hG������������6� �n��P��������{�?1��Gx[$�Z�"Gڃ,�n�}����� KQ����M1'�'<���~�R�#�{�xv:<�+�yX�DTQ_xt���4!�fɵEv
6�?�a�Q�lC�ͥ7��y9�^�c+��5�mn[Hn�y6���h��$�ᘁA�t����D@��0�X�4��a��Pڐ�&�����6� ]u�d��B�	J  �b%R��c�Y���
���}����0v���kihn���d�A���o�N�� XR4��* n|���[�؇�j��d4������h�z��>y�酟���8�J״��v����țmj7� �Ƴ��	?�����0��/#�����*@�b�˴q�	t �E($ uP���N��g_��L�4(N�*��� �}�4����+����X���!���,��G����4Ѝ�u��t% ���o9�ں�&u ֕�3����[̴`uG��Y����-��M�Q7�<�reRU�]��vDQ�[U.}PP��	�]4�+b�G���p�	YǬ�X;�~������vQ������@v_�>e�屁Wts��ós:?vs��q�D+��j}nw(� ��W&����v���W<�W \���W�� k½t�U]�	f�ܾI&o���GjL6�d�<���)	 ��`E�����-�M�/!��|���/~�f�%��9=�*��W����w�x�Ah�	   ` �F���,ta��9�2B
�㸳�����%�)����TV0Tu.�:�
/�vgf{�#��6+��%i�7[<��>�l���O�Omm�_D�q�"�]?��Q\�<T�ٗ��K��kJ����`%���z'$��z����Jԉ������٧�BG�s�#�@�s9-c?���9v��o����+�G�� ���By*KyOJ�Rh:7@Ҏ���y����9m��*�@:7��U�k�?]YPtj�ȍ>U�e������Wu&�J��hy.�����g�2m���v��I�����p��"�������/����D�2��Iߠ���M���?(�S�� �&��WĒh���@��	s    � �-W����: i1�Ď6���Q�xY
�<Nշ�#ml�����H���)X�#�۱o�v/�ZaN����.|U�P4p�w���Z��T�W�:H`�%����^C�0:�f���F��0�8�;6�*&��Hu]�n�!��s��֭�0��J�i�`9V������fM���|�% xr0zn��l�v��O���!�@��Q��fF@F�>�N�l�8y���	��)�Dw�}��G�
D   �ȲUW�C��2������0~G`�D>N��އhmD����\��'{��X���-bs�z�b���Z�~1���Q���㲧�0�i��Ȣ�Y�-�[}���IsG��/5pL��h�6�����O��Q�8���2ڴ+֢��$s�M�"R��;�V�Z=�m�i��%[F�����B �(�[Gr��,���N���~���#B����OW�lT�Ip"P �� O�t~_f[���t�R����Z�w[i�9RK%�nho&<��H���
����2ݣh��b���B�|h�n?�i?���K��v�}x/�ֆi ����$�$l:xj��(4 �.X��U�p1:_ ���޴yh��� h	̲����_ۨ	X����+��9Ẁ��:p��m�Fq���G�:FY�VCr	���x�5@�˘�I�Q�-1�=��Mt�Ԯ���'�>uB�<T�6��9�<�uW�%ö>�s���w�C�.>rP�1���n�c�P��H�������Cq-�Bq ��P�F��_��̢m����L��4kyk�w�Z]���g��$0�ĎiM�k2��̕_�Mm�}�.�1[z�t�����y�3����Y�����S����=�)�д�z��qv{�Oχ���rt�B���s�)����0r  :���]I]}�E�&z��j����y����i�(&j��h/_˲�i�����*�y9R�W�t	�[Y.q���E8g`Ų�èHA��0�#\*LG�f�����L\.Y�hW	��B�پ��rƃ{��z*�w��oO[�{Fd^z�I���qRj~��]&t�4{�������4�����Q�����B�� ih|`�'���t�x�-B�Uac�}�YM���\[��҄?ֻ��H���:M|M�2��AtR��w7������`���v)�Ms>!�}x!���zr��=��q�.6�A+7S]��8�О�C�2l����7���!C�.>p-�&�4I0ri�m�T?�+�9&A���jА(�υ��`1Hk�v��>/=��3��z61�,��r�ҙc���N�l���m��=-�?Dc|�+-�,�5:�xs\�Ů��S�B*���Bb�`2�>afJ+���L4q.	����,K/�p<q�m)q���~L8�a(0���Ϩx�� %/��WH[�v�q��H�э(+��"c?�,]1�H�f;�=��q��2�ka4K�;u���/����4�p޺�����Ej"bڮ�*ᒵpΖ�zb��mP3:ب�M��V<U��5M��|ӄ���\׵�;L���:+
#�Z�]�@خ�B?(��e��3Rc�m��C�W�f>�g��FbG#(~�>+�Er�ؔ�xf?�;lQ`"���X���ȶ�T���<y�b`��x�q��~%]� |@���w���$`G���/�A/j�����Wo��+'��S��nW�A�%�qMYE�>H���\j��X\�6a2�ڲ�jݐŃ=65 �X=�zVº�4��Ƨ���Yώ���iD>�YҴ�TM�UT��
���q��M������!���9A[���h8�+(z3�)��P�f�� ڎ��.O�	��:��u��Q�_�.�͉����?���[�.�:5��~Xql�~\ZV��=�HQ��9H9L.�� �5��P�;w��@��E7s�"t� �L��ټm�d൯�{�����(�5��M�X�v|{�=���-w}�e�y{��g���d�ޒ����r�����d��Z��KWqyY�� �1�D��c�A΁	�  ���%RW�c����Wӓ,Ih6ϖq��~(�u��=#g7)>hKX�3�jy&�;�i�0��f��#7�mh��&�cF_�X�A�8!�����~�����G@]��KZt�7�����bH�Y}�G#ٶy/Z)eQ ɸ�Sݞ3�-Ce��F�pA����܃�j�]�យE޶�_x<'@��P�Q�����qr|�Sw[�����?�}�;�)�AbD��s���m��FTz)�_߈mK�2�=��Y�65�� �n9�BQ�����J��z�}�)}�>�A���@�ҥj$HC7���&�D;���2&���d�L�� ~�c��n����m��L�)[A3q�~��c�-��E���t ��3��b�U�$��q���-�-H�1�b@�@=��D�`�w4���.����w���?J�B#�YT����#�a��x  S�`��������@ׁ	�   � �����,ta�h�V@�G�������lp�-���d��҄��sv�*��O�h�β����H�+�^�(��*��VЫZ�@ u�*,L񽀰xR�s��U��5�F�Y��O�y�N�I�
�i��0t_�H��w��Ʀ���@�3�"gFu�V7:�n^d?V�x���%�s}���ӿ���}/.�p��,�:�Q%�>x�A�
    � �-W���d��ҙ��A����Og��!,�����q�x�T�&�'A�ΫĈi-#�C��d��^Z�V��4��J0v+Q�oE�_�X��  �Ng��B)s�wl���エ�J�:�zPfz=Q�Ҍ��ƅ���7
�ga��W��I�92 �$�
�#"���}��:P�+ˆ�b����Ӑ%WA^�~��r�a��Z��T��v�H����C�()���.\�-�M��A�=�|H6,�ϣ�0����EP�
�������Ĥ!��)jd�C��XJ��鰅:C"���N�-���!��0�(��I�o�v��B�ե����;�z��84�����+
ٳ��vP. �MT�,ܔ �m*&��&(�yl�H�ʽ����Y����;d�Q�����S�J:����M�`:X��Ү⪤���喟}q�     �!����C�ef�,�V�acX��aU%8k���zNTk~F��J)z����:�M7�g�:�U���[ݖ?P-�Z��{�:�\4*�ot�Ӓi�s����\^S�����;v�x�����J�'