c߲U�FL	j-Z��x�\lW��3&*ri}.G��fkXZцe���;��ᒠ�����H��Q�X�o:��'`	vj$N�T�p@�;n��y�"�mr���A���Y*
��!|�-���$�W�0�[�4���)E_Hp���    8!��_���PtP�)�9f� t(p���q�Ln%'^�4Hr-�d+�FR�V(KDa��#���'m�h?���.!/)6�$�ӡz���Н �W*(��-�	�;��Q��^�� ��*��v��:�0�;�)�aA��t�`���G3�h����J�	j��lR �™ݤ �ՃW1���`�!����J�����x`����`Q��]�us�=�Y|\�lZ�_*�/�<�,��	.LZZ��%@�_m�� �&u#�Q��,2A�9  �0��C�-s��)�+O�p�v�g5���=�:�x���Xuxw!d��Z:�S ���P���]0��j��	����l@�����!�h�n�� D�����(,� ��	�T�gGպ����1VF����:�f�h�Uot��$�y�o1@S��`�/Y@b$*�"��V�/�H 8 �%}����b�+)'�[�ɭ���m����P3s��rz��7�����?}�}|~�����m�� /@��*�x.�����Nu���a�*��� !�L���H��}��V�
=�,��nS�W����7���"S�oǮ3[*ܣ|�s���
�����]e�@�rv��Q �0#���. Z�'v~�J��)�u ��e��bp�����U�k���%�|W%&��H����Ytb�E�#UJ���DF�!Q`��o2�+L�X0!�����`4��9�� i`/�Mۇ�z�I���Z���G�m?���@��� � �M�rW��dt,��,.bA�SG�WN�ǁ����c`
�U���G �;LP͍�%()���.G��M�wf!	CW�
��v��ǈ����؀oT�i�Y�jƍ/�#>H�HҬŷi�~��y�1�p p�M���   �Ӏ�UW�C�����K)&E)2l+e|�·���l�*�j!�.��O|�� �����3"��8f&�/YaK��.9�
V�p��,,��%%]}(3,�䳝#���p���d�'�.��>P�)�� @ӧ
1�u|ɾ��ɜR[������� ���hF��w����(��-�8��nK������x��/�n���6����Dl(����2����\ N`@ �5HJ���m��܀4\t�[��K�%�	��Y�Y�	ws<�3v�ᡡ��ћ~�#��s�%̈́����J7�2���V�GY��=��ޅ�}���1H��c�X��g�t�Op8I���ꬹ��������Z�a�>�5����&��rz	j��z{f�N,�m��'C�st��y��Rs1O�*���c�(����g��`�:7�5�_���.���8� i[Y�6\�a���r�#9㶶������&���/ ��R���A
!oZ��5P$������:�U�W�o��:��$��.��~��?*�Ƹ�Yૌ��~#��X��G*�cs��_f�>�uW���@0��?�=�apW(�����0�3��E����]�<�gk5���/�슸wn����