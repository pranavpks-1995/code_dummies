 ���ĈmO��j�G�؋�b��hGt�)��s �<�zo��MDi�Rl�٩*����ٌ����LE�I��uXW_�T������R�pc=H;�e���)-�jo��V�IX��C�� ;�
���Z5Ź��k}yƂ�l Luq�s�'�<�C:��� 	Յ����b����+.��YS�(�)��A&��s�1d6ߦĔ�؟�d!����U�;�R�x�A�bmB�{��[�J�P�����0̛3��LryO�0��;�sz�oF���l�؈�yu�5��@�N^R���Dpߢ.W��s�E971��Is����L\-�X����I�qQ�t��6&:�qd���0�P���})���8�I�c|$�����.܋�cr0�D��|e&"���k���-�?NLN�"ma��\�o����3�g�{*��&�{��7IC���6�����v�&?U���r/n�7V�qCaVL.�!���Ԡ�UGƾ&�ٿ��݄��`+g��t�WS��=/&�����>�;Cu�S0��kr`�Jm�itϑ��x�+
!��S>%���]|�)6��B�0��"��ܱ�0�\����^�l�eȮ:�08֬�;���ѫl(F땮�@0�;#c8������H��v���g����L��@>t�L.�����b��-����y
��[����_�F�X�wC��[E:�ͦI����@�u��cz$��
:�2R��ĿW�i^4/i���z�f���D���^N���� �lYFyb���#Әq!ko��6����$
��y&�S+����ժV��%ܡ�;-�~�,�Ｚ�"��o���S��ް�q���k7
kG�d!:hWQ���2�5d�˲ǋq����M���"�]U��OG��K;����.�ȱŷ1^:P�*b��M���-K	���h��x��#$�W
�8
&�P:����ˬ!��E��A�fy�>��A6)%Y�w�}5Gp�P:��iB�e�l��a��}Le�' �[\�A
�oQa>�D�"�����Zj�\2���>;(g�{�W.��N�:Ւ�6���BiQ�Ai!Y%6��Vi; l'B"9B�8%rK8�V�<���phg��6��+*���`�����4�~0��d���fF۠�Z���-���� w���q���zӱ��%�/��|%5�bTկ꽶�"��XA�@Gm�z!�d����U�+��!�q�Za4��NZ�0��:\Q�Z 0�/�G�����z�y�{��
]w�H���f��2�믂ۂ���U�/�(h�d���l+�8��m�lR���R�5�� e Z{�/�t+KO������i0b�����'����7�m[n����#�^����.wrk�#)��K�g�I��W�GZ��g��Ju�.�d��"p���r4�����(ya;z��?x߱�K!��������tSӻ;01*RQ}�U��n*ݶ��F��;+	��}�2<X&YtӬn���k9���(��8��b�ω]���!�^z��
!��a��Ş����)�+D��: BÝb��mi�Y:��R¨�%tm2ט�O������H��x����pMJ����������23� ����o��!Ӣ�vf*��U]��pl�!`�y�}��y}�ǎpT�\q�Tf��������٥��sMlsB/$�T�x(�JN�f��������t����d ��n�ʧ���!\wυ�4G1��a/j��-�{���Rp�_���~	{�����rMN!�h[���T��D�t���o�Y��>U/[�����P"���(#
-��d���9��ن�Q��0dep��8|S.߿I�瓪�8��C�	���p�AL,.��/�	zPI����a�_