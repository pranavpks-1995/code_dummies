W+�    !��a!dF�2�Ƣ�� 纚�*�.�Y6�<kk����3��)5f�Ȱ��""2>�(�$%y��*�Q����*����Zk�v@����������l��
�\�����&붲��2�驹�_�n/�?��Z�:w[�R����\qb2n  3�~�ڍ�'��F��o��GuuT�    !��=EB9FX��n]Z*! ����@���B���	( �j�F:���ŏ��S��c0�u��/�m%�J�I�+��y���Յ5`Љ�כ/uM��=~�2�w|,�)B�cuZ�w�8�7S�䵿�m��J�&!�!� �r U�i�@�P� ����@	O��1DD��-#wT�II�T�     !���H)Z4�V**��,��ݗ�e2>˥�<U�ȩ�9[�fk冲.���k��c=�w=�_�4r5���n}��T�i ��m�P�>�+�
"Ɨ��8��1�Iˢ����*fؒ�C93��9�;~:�B�7��P���� U\(@@ ,5�>y�_��a�Ɖ��)�
D	[��R ݤ �csZ��  `�!��1��`�� Q�"�$M���H�m:݌��BQ�Y)����9�bwS�� 5���f��[�RG���D��T�����Md#Q�c�����!t|��uB[=���ܛ�/XZ4�>���34!0�M�Ț�Ȓ�BB�pD��o������1�� �gv˅Pgo�Ϧ�_߈ %-�7n�*XK�D  �p�_��   ��0����C��6 ]H��`����{�(π�%-���,�(M5���ʠ�y��.F��8%��Y�]��Tނ )J��w��W��R	��w]�k9;}	5D1m���K�tI�C��B6�j���o<�;�?@��.^'f���1m�g�u�!�B�;���۰����}����/�
������OҢ�R�+�uh��#v����1�ZI�m�y34�;U�P��cxC:|XR�O���k�����N�BU�����C>�~I�k��$�?4A��r�U+|V�A�	Ó�?�5��me�ڪ#9f2�e �п�=,K�&�q��Q�]�^����$�d���fU
M�⌭)� �A�S�	'w���X��]��w��\Cr�p�Q��c��Kc�t��S��r�����qeb�c�},P�����"|�4�Xfڅ��I{	
�!ԛ����L�@���]*�&���t'��5����c�S�Q��m�EO{�bx��L�)�!��"H<�%�qB�Ǎ7��#o�sP�ё��
`ځ�a �@[������4�ȫK��89��1m#�P�NTݜ6�

�1(|����^��!����q&��ŷFz����w��,|��3�,��(p�j6'+>��L|����\�M�'��m�Q}��O�x��L���ϙ�:��Ifđ�j9X�u��δ���t�����|�t�y�4�c0�P�UR��?�$atli�g�À�,?�3� ��~~+'B,v�`@�Bz��<���J?�n�e��O;�e�d�z�NƯ<�H���h-��3�'b�e=b���I;s�)V��U���f���H�u����}a���s�ă=�E� WG]��xg.%8�)���o
���"t��������ͭ�w�\e�����ȡ�2U�]��>|�p�`��� �J(����(ܻqo�7�7^$#_qG�0����Iۢk`� 
�0���IOtP���[��iRC�L,T$l�k��K뀮<J��!9�<ݧ�5
'���`z��D�����5�K�,pc������b��'} �����.��frxs�LIC)}���s��k�kC=�=v�q��>�b�}� ��rN,�l5[�@�V-�a�{+m>�e_����+�M�{Oo�1�jdxl�U��U�� �G3�a��P�]�!��)Ѕ��~��K1m5Z��������+:a��AZ9�Q���?��ib]6!�D�����n�ߧ���x4|����f�aR����M���Z��J��ϾW)F��vl�0��������|T�k1`�|�u/��R����Y}i�Х�7�۔�Bo5)e�$���m���Ū��bد�O����e$��1������w��ݺ�'�Fw��1V�#�m�X�$�����9�ġ�i�Y�]��_G��+����R-+�#�oԫn,`��ʘ�;Ng�LE����2����+���=��<%0������S�e�aN��7 }N��l��S/	'���HZbR�i�K"��C J���[�������Y����Ak������_n���$�%���  Ui$P����<8�ۨ�h6%z��ݣ=#��:����H.�a�(t
�%���	~3�4��o_�V���?t.�5a�2�F�vK���gv�~\X7;�4W!n�/`$�Bc^�T��So؋�V� k�+��p�{a�TTG�ٳX�	ۑ�(�\�P��?��x@Q;x�hfb�c:�K�0����kO%���SKU�P���(6�J�:<0>��.WV[�m���d�Cg�y٣l���NB"�{�� ��l*�l�)e���[�(�c�	v�����A�k_uǐ����hd����d�<�¡� o�2]ʛ D�j�T�Q �����A� >�+x���V��#�s^��iM��iq�><Ɵۖ0u�>jH�̺O$@E=�� ���dȽs+�vP�K;#��z�q@��1o�R��Mx~I2�q_�g��]Rcδ���V����;��=@���1x��/ r��_�t�����þ�[o7��Na�����Tn���O~f��