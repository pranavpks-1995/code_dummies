�\�L�b��-3��ۿ�)�L�c��FE��Oƾm(���[�ZT��{Rٴ:���A��-T3��]9�x2�$�=���h�?�L'�3yGv�+����ʆ4?fl����I5��Ӟ�U3��Q���Y��ּGy�.4Pr&8r�K$sj-&UC�#���4��>P��k׌=��Oa��(��R�Z�n�IT��!²V!�4E2�Y���.D۲q*nd����������)Sd��+��?�[}�p��_^m���Ȯ�_cȼ15����(��5�.�p]����0?!g!ޓ���������/���  "M��U���_�(c����Wo�S��/y�`�t%��c���|V������ �4{˨]߾�ut�U��?jJ�.�p7A�0\TſM�@��Eٜ�R0��{�~Զ���t��+�t�.r?0��;��J���6A��LQ<_�2�9=���D3TQ{��H ~�IRn�窍̰Ei.��sB����+�Vo��k$ê-l����n��&�С*�,����s%�~9�/�PL�~���c�]�2���r,sl��Є�=0����{�5�q��ѥ�[�/Xt�8]EZ6�� IП�y��%V6_x �+q���%6��!y�/\k��I�fQO����1=���\h�+�f �$
��{�c�'�V1|I�H��*vu���g����8�P���'���J9�ׁ`l�q1ZM&(BJ=�-�|�Ϯ6(���0��l���PBHl5kB߸�XLv$��P¼��7O,j�P���u��!�ˡ+Uq��5�C�>>#K 7�s��V}�=�W3H\#u��{�z"g�rSRw�#b@	;� v��?�"}M8v��N���H6���*�f���t��Hm~��S6��T�ˡnh���I+L�@0K���vj(#��a��]����;$�N�8;XV]�Ƽ��*��O�㽤����q�-5k,���B�k��0�:P� ,��?$Oڼ�(aa�hT9�����쯃3���� m] �"�g!�#tM����@�%�!1ʏ��^�C��r:8�R��ьH�VV���ufy��˧�1f�? ORy�˝V��CDL�X��������������f�bj�zf�6c��y�ǜz�2�Jجד�����1�qL����lX=WQ�Db:�X֣k(�)B�7��|T�K1�Bp�Z��Q�J�Z�Z��T-��)|�	<R%�±Z��Z�u�w��st-�aY�R��� ���z��B��&N�D2a{ށP߻��x)��z4$R��O�x[NF�[1l���~�K-�Y�O�A`"�]| [��6�_T��7sSߑl�� o tvj>����[�9ڍ��Hb&��D��A.��	�ת�2^ ��#�MR㘥������`R����UI&L��d
	May(����D}�=)ސ7s4nII�ZȞ����X_9�3�[�8o����NY8y��@11���fP���t�����X��j3��N�`��,r�S�;�,�|���6���{"N��A0� w��*���K,\�(����[H�i���\�O3�Z�_�d|���V�I���?b�ğ>6ې���U����^�]gt+�R����W�*<�{br����ߝ�8c��V�N���Dp��̠�ak�����<	GB�zp�u�¦�|xˎE��m��j�BJ�� �ʇ�6�f��ca�Sޝ+?�Y���eNw?@ƿ8*����O���&�-y��'=�7ϥ �E��&  ��'R��c���H���n�1�Dx����t�mq�bY�����.�O������	������8��c��$�X�$l�h�l&�${��
* ˘Y��\8�F�����������ʊ@m��)��<��ŭ	���5�Dd�!yY�4�/ˏ�!�g��*���{H�وxKD��'���S��D/��߹�V�Y�����&��_&ݰ�l�$��WX�I�&W�ˁ��v��8R(�5!��?���.��K�I,Ӻ����_�(&Pf/ϓ��媫���ԩ��Η�b��o3��J>o�J�`|�����[��r�B���۶~&�t���`���zҽ*O���e(=i�Ew��J���u��8`Q
1�I$�`�Ƣ�7S9���U�>aY$������A;�H��l��Wke��`�d��P�$h�X:^���#��Z��>ژ홿�\"�n�Y̷�w�e��?x�#t^�HY\�E�o�Rq��Le���\�:7�
�e!o��J�\�	_��<30�%vu�P���R�6M�%�S�J�\w��Hv^�K�@�y�Gc;�]�A�,�[K��7���.�c�K"�?螠�U~����E*�����h�?2ڷ�#�C\X�z�ȷ#��}-�����+��������:�abB@�v��)6���1�go��z����X��i:k�1z�&�$o�ţP��b��`�76��=*3�Oje�5���jZ�el��}H+����g�M����2��[~�B��P���ͫ/��9B��6:3�D��i�� �7�k�]�v+����@)}Aq@��_̣��5.���_A�~�B����)��TH����"n�3X){M��Qƅ��@`��)`�x3`ES��
����Y)��F4�b��#a�g�+���
O������O��̳'ڃN[zrv���Z�y|kV�n�5�,Y��2�+����ZWDzGۍ�����1LVO~N�lf�jì��8ءP�1@���j�D��:�>��@mb}�"K;�qWg�Q����k[��+~\�_�U1`�����y����8#�V�
���~#��y�l!�]��%	T��7���0�Vr�sƈ)W���U�+�1�Qǲ�SP�9�a�N���|8Pq_��x��_%�꽃1��uL��mf3����V!�x�U�#m�I�+h����Gp�J`�In�����a� �>�8�ޮ&��SpM����
^���B]S�B~���Ch�Cl���/55�I� �tY{n�EP9��eY��tJu��82f�|��"{�=���sJW+��ؽ7E#AG!]��I�rUK4ɝ�l�ǰ�7O���ޒ���&�?]C?��n*0�%8m6"m��ǐ�2�p�8۞� _��t0ȿ�vA�e|�C���  x �f�U� HX�'.Ax���r+���=�N{p9��Z
��$S�FK�����=��t�V��R�R�@#������)�u�[�I��%�h�
��]�̖2'"�*hf�Δ\��'6)?����9;s�8�)A18�#8�P*�JA�+�>��-͸U�P�ߨvu�p��F �@W����|�,G��́��𛼃�@(W��W����sW|EE�m�*3������QXq��Տ?�XB�0�zΥ ˳�3,
��_s���asL���:�L&���tc�}[���ߴ�uPZi�8�JV�D�r�	��d�]^��r��?B�5��<Ae�����եln��C���ȣ�DM�D��?R�S�<����:�X ��N.N睡fj��5`�f<m`���/�,�~���J3`�Kd{�Ap��%)���ڜ(��Bn�D$(��;�}�Uch��C��p�T��P]�UL����3ZAr����!F��c�nŻ�fa��ঊ�4։�F�ϲ5�b��5���N�!���m��*^ �)|���nM�Thd���԰D*�ϓ^s:?�C���*����!i��
yBw��f<��S�\��I<�sРR߸�#	��WO|ၑ3H>-<��Xl�I�����ٍ��!����B�����>'���5��x����M>yx>F`�\��6��o�Q�:��$٥��8����0Ŗm�b]ͥ��+A������~@�j�,Ԍ�r	�i�~�Sy�]�H?��>L�5�~��n8�-��#�uB��c�L��>Q�ד�>vz��-{�����`��O#�N�/�(�ˣLRxo��Xӽ=� �<��WU�|G��1�݉�>����0.E�N�"'�C؁�   � ���u� d�U3�i,��8��Q���(�m�7�Cr�yR[�GE4�r\SG�.�W
���Z�J����c�;6�rJ�	Z�,�~��bD{Eg�L��P����){ҙ���j@���>��^rH�!�ƞ���@F�o��&�=f�k���[��hpӯ+�]Tdt��}��s;>ؕ6�7JX��[fY	�zB���I�z����c�6kU���E�/a
CN�E�����)�S�_k3)�m�KYv@�#�4Nu�a���J��PWV�m�9x�l��u*��U��0�C�V�u�7�b{����1ulV9+F�z�M���m`!�����ȧ�-����o�p�V�UC�+�H$���=�f�O����`[^���R��G)k��Q�f{i��	F�vh3h��]�D�U�sPi�Hn_�������F��[6�bK��BK��zY�l�Y�ੁm��1�s��!`w����|�IJ�x�!�2�P.?�1+�yj�O.X���w��%d
h�w5�̕����f�Qw�L@ͱ��M�~�z�*3l�i"��>%�Zic�v�[�I���F�(c�a���H�� >��u(�/+�2�Lx��s�\�H�{� �6��=�g��9�<l�J_h�\Bb�MJ��6����b'��- ��2�����aԽ�x���VxH{Q����3�o�[y�k�D���� C&�9x�o�=�\hKz�ŻF3�u�_�����	����:�	�i>�+�s
�]0�%/����� ���a�x�AU���߶+��2R4������ ��B��-��=����!U�24�5g�e����ǳȩiA����܂���ʀ�-��3a�{�ޓ4;���h=�d�a.Θ��~��?C���V�n�����%� ��Q�`茱��y����+�'4��1��%yR����E�17E;�|��$ߦ�vn�B�eͫ�B}�O   u ��-���Ï4��Xj����,7��r��pa@ w�v�$�i7��{�@q9�@���g\�4���Z�P�EՐKZo=6l�s�Ɍ�b^8d6e(_��J�?
���g0�č�AE�_S-ښw+�]��`��ugg����F52��Y��r2�T�K�Z~�ѫ?�ؽ�W ^!$��č !!/����^ŕ��+(1��5Zؔ�Lx��z{,���o�-U��d0�a��������~��{�Q�s%���W���Wy�̤�����V���������z�b@�+��$�[ʕ�u�)��bf����_-t��XK��
<���{{��~�U��Ny�t�4
|D��ع���/,j����lF0�*�EX�7��� ���R�j�l���P��v�qU�tCz�>欿�!�ڋ>��)�~�"�����!�d�Ɨ��vM�Z=e�m�HQ��v����F����yf�7�u,$uO��r�����3�\������lђ)� Z�c�*�(���sl�`z@v�ǌ�x>`Ǹ��+7���.	������Iq}���ANv�T���@��<�F��ÜDU�0�C'��+$.�8N�'��xF�+(G4�{�è����"�\]���� ��M
P�T��	    ��X�U��C��]0.��qHڮ�A*����	C_%��F�(���*#�<ZY�-g-M	�>���H�z��H�h�Zx_"�;�R��ś�Q�ª�<8���V���9�;2}g��W�=U�n9�r'�TK�uV��ٺy�&�㾯�	_��oo�E�{����r�x�x7B�Z��G=-8��i������w�o���c�cJw�����	�(p���#;℗�G��ŭ��l
�,�UG'8Q�~�s�C~хF�x|�1UK*z�4���G��*`�'�(yB�9!�f�_�V3�A
o����,_x6%��{�;��rV#*��=��ξ
mxh�A�M5�c�f�[��F�Z�5X�Y�mZ�ǀfx`��B��<�'cw�Ky�MT���B�Ր.oS) &�~g������b��e<m�b�͚m��Xa�]���Z�SR	&�K���7����'�+IWB�j%�!�)l��$�弶��	M��\����:���� ė��n5V/Y�:Pwn8h��L5ψu �kL��2@��10���*>�1�s�p���i�Hk��4�J 9��:㪷��:�A)�:���S�Yf#�u
��(�PJ�Q�`������o�<����;���d����ҳ�H�.(��<�W�K:KV~ۅ��27�Pm!\���Փҭ�&�o2/2��i�|���r�!����ުHP`�e1����������/"QrH!�C��B3����'��L^Dέ�)��]�	�����i3G�m�qE�43��K�ʹ=s��M�l�3���r���}A�%�� C�jE3�À�n�c����i��3��%Z�b�;A��Hqq.��CB���v�3J�Z������󔔪<vg�t�渦��34M���-9oy��k�P�!�Y]^�G!hb�pћ2��g�c�,���?����ImɎI��)9]�$�v3-��<V?r�ix���и(����xa�D�X�w4_u&O���/I�z����������ԣщj���8���ɣ>��SL�Ke� �VH�a-����۲Wm:$�PM�-@vB��ȵc�ޓ��D�W�y������|���"��\�ԕ����m��ˬ���%��BO����-�����*�b�0�+�����[�F"�Q�a��1�4ѐ�do~G
$�����Fؔh�+$��{tβӼ������?5?�$BVW��u�ѐ�4~Z�觉*�90fq�h��T"�к�f\'�ں��|`�