p���kM�ʋ��9g<-C%���$�r�w���D*��]��5�^(��J���x�&J�O�6u�~NG)*�E��!�zbe��
��t�D��n���+y��؇#b�M�Docr���ی���%��7�ݫ�1�ݓ�s�@��T�=�,��(A�;�
=H�ɼ�gJ �j8zR��T�D��fl������U��vhC����V0h�b����f3_��%ŝD���^Nx2�>c��]/������kٶQN'{d0��Ԅ����xSD'��ET��a�y��J�.F���o��-+�r2,��^�	�eY��f1�pE��=LV���p;mD���K�!�����3;�G�A��9��;}։�A<�?J�BGF�c��}ϗ��1ky洛.�jm��q ��a��.1�m�+��zm�5�raP �U��L�U��?��C4k���OQ(;��ky_�iQ�!���(&Ԟ��2[�
6R��pm�rÝ�Z! ˨�;�=:aa֔��$G�J������v���%�|6�S͝��<��~���o��r;QJyXuJ$0�Ѥ��]�\؇&=��������z��y�i/�㢀Q�%hX�$���	�/'�:�r ڧKmB��7�wC<g9��n��1޼�db���pS�"Y��u��kpMb}-�B`@&(:��B�6��(������2_u��՞zz]lQj;��̺���yw<���q/bi���4T@��:;s��Mΐ��0|L�RV��'����Ԩ<�QNY��z�;�����M~2�ڗ7GKu#[<� ����|<�~����&'�8�B�wFќ�sZ~�[�6��#l5�����6��E]�����6^gl�&J �xf����n[�#���Q�Q喃�n�*"��_�`���'ًq&� r
�� �g���,A-B���	yK)R]��iw�!nW�>��Q��ΘM���-��_�ӹ���6�Ȏ)�+I)c� �0�!F��-�N@����q�!K3� �=Z��} I����_!��3�ϴ1��֯=���1�V:ZK"��|�ޱH������ ��$s�/�KZ�Q&����!�ݢ�� 싕���