�g��jQ�v�BC���bʚ�ʖ!�:�������U�H`�5W05�� J�vݤ֘��v=��%	���LW#щ�-���/�O�9S�ɯ
������f'<���(	��g����*��g)��H���FBL���DB�X�� ;��N��wnJ�@�J�q�>��Hb�r-�QbV�G��UUdz
hj�#mW�^*cJ�0��º�M���F�<�<H�J(߰�|Yʻ��k];ϛ�����o�%�v�U8&���|ײ���L`�.�òy4�ŸB��؍(:���?`5��k=A�*���&&�q��A'��j�&�<Œ6���7fQzR6z��|�CO1r���-��	ӄ*���$��}��ݜ��Z@�z��
��#z�ڤ����&p�lK{_6�fs����"��%ʦ��ĳ�VԀS�Ħi�K+j�W�5��f�}��&��[��p���c���<ٰ'��4�Ű����8%����C�^�"�5���϶E�pL�v5h�]�O���Vؼ�i��a��h�ﮍ7���vcqNW�
3�Z�_��>̩�F���` ����Ve���Ց��)S,T�����c]��U8��]�]S��]�� O!���<���l4W��@�[ C_����"�d�G)𱂯�gH@Z'��� ���S��
��hu�}�?6b�#"�~�8��/$�WC���^�p�P%U�|�a0�[n�ay���3��ψ������{��a�	r��zs8�: ��Z�����RA��O��=���7\�i@;��Q���ǈ�1�iޠ�����6�U#�����V8����}���hJ�27�N��hR]̀�/�_��@>�<	� 	 Q7<�|f��I;��s~�ʍ5ɚ{�\����ZD%�`�y)���Z��t����h," ��LHo�^��h��� ��n~�~�	r�KSՂ�j��v��k��r_a)��+-�I�Q3�3=R�2�T$-�ąrw��no�PN������a�Y�7@���:���b�ue��9�+��