{0��j�����f�C���l��6q���5�8)He���:��2�/a������^0W��if7%y�i��������	؆�*�?�;��J"�l�WBioF2X�&{z�f>�ޮ~��#ޑ��8Y|ǋ� "�����Yh++ꊴzs�[1 ����	�7҃!oS�z�9�󈃞�!���-��@�Y3��s�t�g�Q�W!3I�-V}.^z��i�Mt�ٵ*�@�z�~�#�q�`��s��6�{KG�-����I
�}��Zl�	�y�g�+�_D���}��76ׂN@YĀ�DK�f  C�b'RW�c�
��5�8-)6��@��cvk��r�pc���$��� 
�,�!D��DaN�F��zpK�\�S�(��(6��˓����^͛�A�q��t�(ШVs��X�l챖��Q˘��`whj��n�qq�2��YW�R�d���<�{&[����� �ݩ�����WǑ����{u��Έ��6ζ�-��O�7y����XJgл�m���d6��m:��C�����ي��=�o����0m�ԧ���ˊ��
�(��x�u�GP�[6o������9�Te�eC\Ѷi2�ӬyV�!���ДF�Y-і�bd�Dm0�<Qé��оox+�a)R�m�kX����{#Ϙ]mE�i)<%���OM��F	>�W�q���MD}_���g?�%���)�wI�vEcg�Q2�h��>��e(�u���0:@�U�|����z��E�\��E(S�Չ����o���&�����ż?@��n�c2�@h�����3u<c+'�w���=�xc���� �٢@{"nMrhT�18�b�˅����a��JK�������6�M�:j�hd2յ�i`Ȕӹ�]Ϧ��׋E��W�q�_%�%��йȳ&��*�7�k�\Ӱ�;켦���"^+z�\J^,�[���&,=
��)F.���-v�� ���?�|U��4:X�|�b����>y0�A��p�e�8kT���7���#��ji���~vIT[�zԺr���)M��=����xs��;Ǫߧ�Gw�P��x2�<�&��6�Я���?�	4��q9g _�D�1�C������J	�Oْ����-}��S�hV��ީlv0g	%`8�G�����-2����1��c�X��3�&5��r+��]��
,���M�������0)��Pi���#nRnr[t�'���|�æ���'������)���v�'}m�w��
��n4��nX���:��~�-�될V��@0_�z��!V2��	I𣬙��+���v�ރv�1ߢNW �1K�%A��`)Y��"&M�UG��"�/q�& �i-�>vG�<�uk/�S��������/����CJ�  B �&�U�r����}W����d�E?Ѭs�0�8䤦t� �ۗY�ǎb�&� t�M������+�E��땢�^�#���Ċ	L�U�84�gC ����_y�Ʉ����N"u� P:�
����'� .���$�2y#�U���` �w\.��3�}WQ���v,��ﲋ�M���� l�����"���@��Jx��{�D�CNq}��� ���䭉�݈�j�`��O
BӠ۸5p언(�V�Cr�"�ڪt�1=b,���g�G�˟�yW�Bs,�гd��:t0� .�!_I/��HT��q���'�f;H�A0z)Z��j�~���
���EdU"��&��VL��`,)�Q�g $H*?���4�6��Y)�s�G�u�@�~1j�eɂA-�`�o��q\:�ȍ$�R��k��%�L��i<���Oݠ=�f���8��x�m;�G�꺴�t�Q��%e7}3ݺ�~d;	�z��#�hD��^�7�QI��@܂�Rv(,VS-:v�^n>tI�Z�K
�)9s���.�r��v�ǔ������{��]����EӪ�j�iX&;~�I��������3��g4�k�c˒�㸩����EvW�V�����@| 4�U;�n���ʜ�C��V�^�ۦ�����N4HA�H��K��o����l�H�vp"8�f!R�T���O��^��ȇ��(3b>��C���oyu��K�l*�YV���V_c�N.�Zs��Yn=�cC�y:�ڭ䀅�}�#�#5(��{�PT��vS "��[�>�yݢ�Z�t3ۦ����IH-�gL�C9�<   1 �F�u�sD�9�2%q�@��l��vPsS`ÞzH Z��6���B�(7�j#�A�Sh
�e$���x;�.�j1�2�$(����������b�W�Z�;Ҩb-�T��L�u};��Bj���]�S��!�������p�g:D�����%�tF�~o�%f���~�e���ƠLǁ�������I��G�aKͯ�ʴiL����{�>�>R�;$I���w�'��T���Z�K'@.P$