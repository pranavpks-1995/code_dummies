�bP� 1��>��A,򭯶{H\<v��L��[��u:��1�]%��-���\�l�.�#����mK�������oŁ��Mz�l&�6�2W�W����*f몎��x5���8q&��f���y��ol��]�?ZN������sc�m��:E����\�2���z����h}���j鱦�V�HL���qF�^.�k=� �i�͒χ�4tl"�K��`�Cť��Ba2L1�V�ӭv�P��1>������c)�LP�L�$I(��UNK�矽Q�$��it'u1��)t	w�3�p���{��{"2��!���z�M��+�[ݴ�4����4sM��LS*.��n�Ok�F ����B���ә�Ɩezg���Z��S�<,oя���y\ �,8�E��u;n4�
*u+��8E|�x�����f�`�)�C۪�1m5�b�t�Z�z�>A~xM_wܚ�������_�8�r�sL��G�I!	���\'���J����:�ڱ�%��/	�L�3Һ����R^TFK�����Dk��4���h�-�w%DX���e���� ꪏU��e���MǾi�%/�X{��Z�힂�z�S]����']T3$���Ѱ8sm��Y���S�����[�.�l��\��:}y��e��(��>~�q��s}�̣T��Ʌ�z�!����+�?���` �o��O�4�Qsp��*rR��X�J�ٵ�N��MR��V��G��~V���`��gaA��	�I�Ц�&�G�����HnI�"Z�����gt�c�pm�\_h�Օ��Z7�CcK�t�0
M��8c���O�l��N���g&J�M]��`Re}�����L1O��:K^%�람�\�S�mU�3#BX�%	����N�k�����)K#.b�2���u�
$	�՛OG��)I|�\zñ=_�m�!����ڈ�ʛժ�@V��3yLoM��r�Q�.f�nsE�����/���qc��Jr)����Rb���Ҧ