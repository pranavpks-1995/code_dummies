�L�"��n���['?���)R'^��课����h���h��W���h,��n��x���	���J���u5�zHn�0M~d��3`�)�@fl�6�W�2J�t��+��ev�o���Ի%`l��C��ڣ��$�\���do����^A��7�X��?��`��"w#|�$�U�Åq.!io���t+��،��M������;C�ޟ�mT(Q:5�zI>7���VR�U�Q��M����?B%:A]�6�l�ʀ
�ך^w���[�4�*�5?����Q�� ����ګ��{�{F��={��& � $N|g,� A6L�n���8�Ƥ&�5��&i� ��x�]��!�cs�X䭩���z�w"PN�]���<�Wat0� ;z������[s�����7܅Zȃ Ɯ'g�� �d��C���T���T g��@�5�^20��Hh�:��u^��Aːo���-��Gg��8��E&�!��������!��-w5M��ζ��@<<<U���;�bګ�Ѐ�/(ᥒŧ�7�AM�WE��3���9ĥ��u��-tiV�h���RL�/�5E� b�G��� tU��rƳ'�a��7�"]�������߰
��{�KE5^s� כ)ƹ{�$��!R6�ܶy��hZ0!� 	����= ��^�P�[��Z�.����,"����ȅ׊D*������;�J��ȕB�$�P���8��&/I�X� ���r���/-�`�m<�v:�m�л��|�H�ȇN����2~�b<������
�	�8F�ѺqMz��HUT&2�m�`Y !�葊K9�[l�@=��{4���2a��iuޟ���O�g�V�r���]z�iE�>��DD�h�[U��|(%e�&�,N(�P�,��D �}� >�{.���d��`���D%>��?ox*҈�Z�\DƮ�1v��8c��u�[L���6i����1��( p!� �8 Xa��.Tc�~D�	�u�_6�l?;���zn68ŖUW|ܭ/8�8�d�Z�$n��׼ �# \����7��@�r�@��v>�>�� vPN"bu�4�8� ;<�$3�`�)@*ػ4ڢ*SxF��UK��m�Z���'q�~��@!�84�f����c\Xΰ��e���Q�\���Pak=��$�����D F��-(�՞֐* ��;\9  �*�kփ��I���~�L�_���Ru�$	(Eu`�o�1LI�X�M5�D����o��C�^�����R�� 8!� tQ�}6ƕ�h�Y�������跘��+�_��Y���T�A,�O��k�ӮZ��2FӆM�8���UX\	F�U�X�p	��ð}6��$����J���cnH���W�G���&�4N��P�m� �-�*-d/�T�,#9�$o�U�壜@l�Z� �!��X^?ua�V*���6SN8{��o+���1l3IH%i�>�ab��e<���U��4)1'�AB��Q�����F�>eJ<nqAA�'A��"D\����7&�3��z�o@0�WT�1 M;����Ӭ��X��@On���Qe��h1` !�r\^���+ |��p�u���D4E}I������o�U���w�^YM��Xĉ��Jަ��m��":(HIi��D,(��$�(@B@���@.�Da:gY��)���O�/�H���<ȆQ���s���>����!uQ�S-� �P-��   %Ұ�UW�D:0\XV����a�*�0���Z\�,Պ捝[�=�L�JBM��ASv�v���;�L��"�g�ǜ�*�
&{�R7��lR\L�]�s7�ytd�C��?h��<݌�@�ABl=b�Z^��� ^�	ڠuag9oY-Y�s9y33��1��Ŝv����m�l��r/P��}\�V�q�5�X��v�F ��M���_���%�z .��fHt.��0��u�q�{�$	(��<�y�6�Mx0G�5�~Ѓv+�~�g��(�jV�[n������ ���ns3}�/B2[1=�S�H�n�/��چ��7��&g�Z�u���l�
�&�F�şBGMS
���[�ֱ�o�	�с �U��Gs�V,�n�IdA��l��g���pċ�>