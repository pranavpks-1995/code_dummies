��,h.?E�d��h�:R�_��o���:��_��HP�|V<{�H漃w��m��Y�)���r��#EQ��L_;7��L�4�Z.r�D�b��-���2��(�%��X�sp�R��mRV�dSK�1[�#>����?3�I�:l�+n_:;���c5V��J���t��L���ŷ���+��x�V�(��?�^k��Ԩ��Gw#���#N�P$���ek����"�p;�J�$I�0���[�F�U{OT�y��㳓R�]oZw�u�q5���+��Q�h���hʳi�5'�[���+�F^ 
�8/�P����-,�B	��V}�W>�9��<�ޓ�Dl����Lʂ��h�7h&�^O�P3�EH�ʂ�������!��xP��o[�h�,@+���{Ef����x��7��{j�v���I_gf���}Ѱ�S��
^O��GaD�g��?ч�8?A��S��gՃU�5g�~��n�i��ٷW���	�Z� M1����dk�f+k��}�F��K���uj��@    !��I"B�P��
P �h  �b�_^���`��_E"����W�4`BU�4>w�B|��F�c�H��߿1A��o$gf�-ޒA��S;���_˂�teC��� �la暺�MG0�}S#�+ ��<߰	�H� {��朔���7uPIqS6͔ 0     �!��4ڋ�n;2 #�'�����zatN�(��x��~����م���P�%Xs�l�hw����~�)a�|"�nKrarп��=2�K�I�A^��1�6H�{������(N�_N0<�i�i(S{����TbT����     8!�#1#A/*`CaQZZ�, d�v����;*!I����p��.��f/���#x�yq�2K�3����躋ֺ	*F��aN(R� g�����Sa6|�L���s���T'9  ������MGʼ�鍻�;�#8��m�
K>� dˇ&Ae3���=#wU-[�s�
� `    !��9�B	�Yb�A�B�
��EU�CE1�����|[�R����/�X Ɛ�9�4��Vr�D��ȉJ 2*�(��ۊX����{�K:�|�����P.��x$��Y��\���@� H��� t&���(q�NJ���0&Q�4B����Be�	\�H��F*�(|�T�    !��UES) ,Ph �ة�i3S2�t�L�J��M3fP�#dX�0���\�V���U�kͻ���\��+e1[;��čP��ԓJ�g�$p�7��1�s}�	�BO�S7
=1�	�`$�	��`(�����\s��tKp�a�ͺB
�bmr 0@�!��X�E0�ǎ	��- ���&�� �)&S�FeF��VkՄ�Ŝ$!j���2�&�	:ӠK�ڜR�9��"���z��K��Oj]��*�J����.�&(�J�4��@.���j�>����Ϧi	 ��`�9,p7��]��G��(*�=��Z�٤*��%V�`  �!����$�yRX � I��(�)��ҹ��=�H����k4�,!dϱü�t�6�`e��A�1Nk�����z; 9�
B��a���v�@x%i���Cv�"�R�6��A`vp�'p�oȸ{����'�O�:����m� #UT�$v�J��@    �T��   ��зU��0��N��}�3S��9o�mF��WEm�����x�����rw���xS���������`M��1�"��ü��w�]tI�[�]g6�H�P[]~8]�����I��
%tZ�dJ�E}��E��)Ⴗq�7zF�w��&[���Vu���[2�Y"��I>�v�X��T�s����v�e+UЏ[���_5�	�s�
4=L���`��w���$�>�>���?��}�?9��Q�C�O���l�!e��Ú����:�z���(���Q��KO��Xa�E)��� 13F�:���I�yy��H��#�ӽd��v,�)Yb���lt�UgMX���D���B�zP���9����WS�r���Ҳ(,.3��v�[�̳�A�7.
W�2RYH�.dsr^e�M�#G4m���<9 Z��c܀�B��V�ODr�T��|/���G��\v�-�ĺ\�<bI;D{_����gp#�BϚn�]��|�wqj�~bX�H�����@�p�� �Mw��T#1�T��dUa�"��a�y<�*ɒ�;1c���3M�o�<2�YPx�(�s`(�`��0C��wޡЋlvN<��M?�$��?kd�M髂��9��YA��-��9>NC�U�k�ew�~
������C8p�Y	U�~āQd/�iX%<��b(����%�>�1ݛ�p�Nc�������c �ڏ=��pC躁��u4+�&rr��8I ��r����qTE�HF�z��� ��	���������Za]jH/��SZbŘ�|��"qS��S���UB�H�7��v���H���++�gg��^w�/L��������4��B��E�����Rf����ܽ�+��b5���1�z��R�ַ&կߎ䮐�XK��U[}#/'�e>kq�>���)EB<�b�5/0���hC����0}���$r>���~`��b�N�l�G�:��޿£&/��~�(���=,N�}�:�
�B����)'W����m��-�(���#4��x���*������Kz��/�֫a�f�Ļ:|��c��Uȷ9q�D3�/C��\�N�:���`J��bG ���|����W����L����@?�6ohb/2*	���� ���@�p��k-/V\��9���}�L[�)�T�&_Љ�SX_O~v��v�!��D%�mv�Zrt���>��������Y�����%�-F�o�|ֺgý�0$�|��!�*PaT��J���#�68&�W�v�*]in9���G��9�Eʿ����=�{<����w�:&�l��렯+d{v[�	b��@餔V�.�p��)��>,��,�-v��Z�E���_�-+^��հT��9��mO<�����
�i/Fު_[?�-]E���
&>r���[.�働=$վ�-b+~~���4�;������u�ޥ|~��R#�OlP�&�c�	J���i��5��V=ӵ\H�L���e��%����ɗ����`��M�b<u��?) L|pQ9�9h�=섎��4�z�O�n)�`��ufV�D(Յ3m#�:��h�� ���C���hv�F�����,���2�T+zmE2g�˗9�	/-�f���QZ�$�z;�Y>�\p	_�5+LXƶed3þ
0-s�d-����`�H"��X��wN�^���4 �����7�A��AK��[0)<�WDԤ�|��Ng�����q]{h��k7y��Y'�W�d��^ʽ�,���wt���»��a҉�1ʡ���b��B6َ+m���ߞ�Tfض�Q��5��w$���9���j����p�	|Bه�c�.D?�wp��PY/�_T�����,��4��,,T?��Gw���;�7eÓ��^ ���Yf�*΅i59+2$,WJ���jx.oh�V��A$H*=�����A&��%�K���Z`�mt�yqSjΩ�>�JG�,~�)o����*���	'B�.LQZ+o�#u(<�W���Zy�:�;3�N |f�͋�U��aOr�4�N�ڜٰ0�����l���8�PV�3Å"�c4��+-V�^B=>g�ybV
p���1��G~��v��F!oy�e8�<��|��C8�1��;�B���9f
SТ����:�Z�*U-ڃ[g�>E�N(,'�w��K�;�=%:g�L�B2P�J��i�Y�Z�[f�-�̤+^�#Ơ�߀�)���\-�ҷ��A��(󀥱�˄Qbd���	��*��.�EGD+4=T	g����i{(�$m]l�nGN��W/[*��eV�,c��� ��=�E{������j��i�&�$*tV�tu�n����#e�V���_�=�z���q��
� }G�� %m���։V���y=�*�q_��7����{ga��g]�٤�2�M~���vڤ|嫈���)�dՉI�	λQ�g���Cg�O�/������	����,�������P(�d�$*�H�me�(�/��)э��Y%�ؐ.ӷtz5h!���/��=&C�g�����8������|�S�:�������ӛ	��x�qӏ�B(hg��� c�GY/?6Mˋ�z'�B�n�6"Ͷ�/��u����,���&TU1>  ֓�T]��Ef��kJ�&!༆e=^��?HG(�m؞��:y0զݓ-���!����PtQ!�J���m2�zr���J�6��O/�"���9�+���j�Ǳؑ(}�=�sHD�v�v6�	h�&���;��izŘO"�$@�1�-�y��ަ�Ѣ�BSos'+$93�л7�˒�ĉ�4?��X�!���� N�`{�T�% ����)��X{Ln�ֈ �F���s�T�%�&�a���
�&����˪L`�J�O���е�	�G{�nO#��R%��	��%M�F���.��B��4��|��t~I�tY/�fM;���a��xD�K2σ��	"�j��ڼȗ�Y=��&=���T[�b�Kd��U�d��<!�K���o/2v��yt~��J�,��^�ΠnE�m�Ё4q>ܐ�(���7cX�2j�4��cR�u�_Y?Z#���,M�|�$ H�����;qqr��,�Kv.'~�6K��r<j3m�!g��M�N��n{�����em~N���{����(�=Ş�?l�_����jd��J�z��맻!W~յJ�,q.q��V��*V������J��8k|a�9����O|&"nRD��xO,L"����V�Q���-���)1nC����^�|�*�2Ȉ�z�݆��ި��j1Z��g�}����������o�g "�N�u�z<��2���?K7����&D�dX)�ۯ��0�#�CLL�?k:���p�Y�L[�����C`D4\���xU� !�#���ju�)Lt�|?/I�s�7h�U@}U˨_M%�B�u�	W��p�+���D�p\�Jua)�|s���j�cQ�q�Է�