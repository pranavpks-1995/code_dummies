ϭ�=��ZZ�+F��w酠�KF�៦�o
�N��fJE��nvíGc�zۡ�Ifo�u�5zך� ?_N]�[X�5u�Q��(�`�\��o�>����뷳�7C�j�x�öv�`�jPO�dLז>��rWv�&5r3���tG�%�uW�^1��co����Cl�?)���_x~�n [4��^��;�s���8.F��[1yjs��)�~��4�1��p�x|ٹs�ij��HR��v�n�
�ՠx��yU�W������	Z6O�Q���Ģ��N�ΒBN�����?��aM�����zҞ�g�e���{cj��O*-��m�:� �V*+VY5�:7�N�FǈBөˡ�*0� �姞l7���p���ܹ+R��RIl��BȜ�C��6�r<� �y�v�a����f��w��<�Y��n�BA
Ӽw�13���ڡ���_�9�v����Y������J�S=G��QLSN���k2-��Hg�>�a�!���^/���9�4�TFs��s��n�̕����j����0ة�p���A�KH��Værﵗ��/�?���)�_��\a�>���*@�0���x�k���چ���� d���f;���*\�X�\f���ce����e��ট�����%�x�44T���ɐ�[ª��N����Q�=�?�[�u�=Y�j�2���sg�:�K�>���CP�7D:;[����-��3�;�
��?w3�2dI�e�vuHu��؛��(F�5k�A3�#m� $��-;U�K��ù�m����w�4�;�u��-�|�/�<joR�����})p7a��S����g�*��y��V�S+״�(�y܂���'��N�+V�x ��8�1�`Y�݀�A	*�s��`�A�p��NY����rI���Cn�B�Q����W�9?�b^�a6��M���	L����7#4��Ģ��H��Q��OTT���1���hN�j�DK"�˦��q^�Q��&�6�w��!��X[�%�\Z	�:X��e�-��j8��Ό\��U�?QhB��a���_�G#�]�9��$w��ْ�ôw�B������"ᬀ������c/����c��K�Z��D���e��޲��Y�n�Xa���w�J�o�Ƅ��X嵟�i��Ҭ"0�8���j��a�R�vf����ѭ�u�gh��S�����h?�Fv��k:��%��_.��|g�v���rj��l���������8��C֘�u .�ųd�����?�Æ�,�1��?I�j�x!ZY)���6]�EvH �J�,c����]gXgE����>��rLm��'ZQ��tn��`�l*��N�SwY��4��d�l�&hhj�f"H�G�ui��.����2)Y�"gtz���H�e��,�`V��F����@�?a�.� ��~1���ju����+0�'u������Du��J��SWܸ;\���E �v۩d�2.�h�HjL����+g���7�jR��ū4�����j�q�'� L�hB �v��e���[ڞu�,n���T~�'��F}�G� \k��V�<f�|3,�vIeu� V���k��r�I��#��� p�!Z
��\��.,��|P�t�F'��\]�H�-}�c0���A#y�h$����V��#��SRi,QP�n�]��Q����l�2���Y�F����8�J6�^vg��!3��� �u�šK���;>+��(⁡Ī=w�՗���C��jI	�P�|�<07��(As��.L�הf���&a��R�K��{P�SZ�(��F6����W]!8%Mq �,�];M�lHf׹$c���-(MWdЃs��λ$C�c��E3
�t�]=
�V��k�Ed�=<KR�S���冬Lځ+	$�B�:1����,�K�.J!&N-0���[��$"U1��?��P����~x����Ya�X�=��(U#�d����@�3��Y
c����^p�#Q5ă��_�Ϥ	٘�J�ҥ���X!� nC��)�F����V�2_s;�����؃fopc	���' �Ͷ�]��cf���ͽ��+��Vrg��p�#����_F�g2�}/z�3$V���kmk�Ҳ�{���˙I�qHM\�q�	p�$�z&�,ap�J����O�FG.�Z�G�@�`mJ���"�$�1��K�
~&�a�)�����N�wml(�G��R7���J'���_?�
kL����wyV��8��r�����"�!I����1�e��V�M>�:��R��}�7Ǣy/d D�O
F��a�����r��N��@����C�*�~��r圆N��M��e�dM#t-��$�����-��[�c�c?դmO�1�[j۔��e���4P������YA��|X���Ɏm��ۻ��k$u�
�������.D*^({|?��j���:�� �8����Mc��E�JA N�<�l�?�٘t�D�JGP����EL���	�5�Y�S6 /<�|%�F�X�7�$D��$"T]רa�|� I7F�J9;+���0)��@f�0��um�O���y���%ĺ?1H��C�� �����1D%��I�%q��.[�*w�ϸԽ�������k}���ٯײ��������s���m��D���L�A�ܔ/&�w^qS���W�21G�+[����*�����
?�����j��$�.��2�]�r�B�%L=���m��xK�mC�&��K�O0����!�1�V9V��Μ$������Gf�F�-�H��-
�Y�H�4�0�g��{��
Z������P�����- �E�W4[0���R��z�B	0K�u̐��Ώ3���~}Ψps�6�Z�T2�˻%���/%�z&}_�F��#�|�������@a~BC��ca[���J&��4aY�66e�A#I�����Gu%k�7���m��p'~D�9�u]n��+�b���
�%v (��es�����%�eO1d�"���i��g4hL�4��=o������3�'��A֩A�V�Ҁc]�h:n�=��O���"�{��7��Q� �t[��O+��lY#k�I[��(Z3׺�:�x	l�٦���w�+CA��p���:����"����͎�J�� }  
��D�xc�(�?d���GKR	P&��^�'�'W{�O�=I�fP��/+�4=E�θ��
"ܜ"���� �6�C�h����s�%<Cw��7I<�Q��	,�7[�@g���옪��p�`v�@CvG�~EÜ�7Y7\�u�i�?�]P�'���(2��^��H%A����]����Xy�V�����n�+����VN������b&ߛ(�֤k9B�Wp�K��! �Z�XٌfN`�V���X��>��v%��l�vs��OH�y���W�M�d<�eCe��2J霤,�(-繘:��������W[w���c~�_xߪK���+(n�6u6!.u*4m'�Ҽ<"Bp2�X˯�I���h�A��i�b�=p�b����(��D�[�v����|�e���H��b�Zlȇ~@�:T��9Esu���,1 �Ce�я'Q�hЍ'=3t��Q�^qa�p�<62Z�u2��bO�5�3�A�J���'(n<��L��0!ԗ�m�^�l��)U�dY���ac�*�#u�n�p�~qIQ�_�md��+(�A�g;����$p��62��O��0��8�t`�XJ.��+^O�@l�\��X>:�ϽT�LlDa+S�;O�=�]��mQ��&�������Q#V�?X�9/X��rT���K�`{4�}��ߡR��p#)����e�o�>1C)�c�R��J,������A����lM.��;[.m�]�$r+�sxe'�?�A~t���������N��	nI:�akgV��z�TB�oD�l��?�?�4u٘9�.���&+D"��a&%.�M��+@o��oRf��D;x��Aa��(k�ߣ��z �����;_�GH��i�iX�9nQ���1E�k�ݎ�Ͼ�
x��#6-�s��E���]��KdM���s���}D�R�V}P��	g/����Q�n�3���&�v�w��Y���O�8;����WG�З�J��t�7��w�p��9�
�jv+�6M��x@��x�C���X���c��7	�dd�R�-Z	��x�2v��UO~�u.�⫤JIjB����4@a,;��^N�kґeߏ���HT��[���9�zT��+�|��.��o�"fW������<Ư�GG�n4����_�	��6��� �딈����r4D��v
�~ɕ]�����~Q��_0�v�r83�E����
|�55���ܑ:��"L�%��rd��ny
�.0j�'�Vm��s+��<*"t͛���8y䶶�gr��x��������~��^(�U��w�=�E-�4��׼�����H��AkB���ɫɹ����@���ShB��x$�	�6�"��*]`�(�Ws���e����,�^�?Өh
�[fd_�~�<� *�Ů�<�$�T���\�O!�hW��i#7�+C���[	(���5GdԈѢvfZ~�D>���z%]�H lVv����כ�&�����G8�i}I�f��L����>c��/p����uD�;1�����0E3����;�X��i�3ֳ�z�D�tF�����M�����N�j
D�t2k�S2�R��kJ4�d�W�ZC�R���D���:��DY�៻XRnfd_�87:���+�h�$����a#��0Hx��L��ⵢ�T>/�]E@�cNR@+��n%c�
	�dM���f�"�ӢS�M	���0�,��2�2�,�%]�?q����w1T�B�lU+�_*t�Z�����v)�>ng$j�k��q
i�&��+]t'��O۵�D"�v���E;Py�W+Uh���o{1�Wo	5�H�"�P}]�Ryih���(%�<����{����=�D����Z+��zv���*"��].E�tA�V�,wK��p��8���C:KyA�'�(�F����M�O��<A5�S�nj�ȉ���t³g�`�W;d��Q>*�W�镯��6B��[.U����7�(��;��%M�N���*�s��O�t����U8�����&��1R��ˠE4�a�Sq~m�{��LQ���hh���N9���K��x�zF�>bj&���a��PÙ���v��B.�r��$�{�����Z�����³���l�N�hp|NF����H�`Z��D�����I_*qؠ�Or�g���6����F��on��8�y��7j�R]�?��~|�t}� wQ_�&�`�ܮ�G�B:ժ2��
�+B��/�I�Y������y��8֛-�[eFѶX|�rKؓ��֌�j��Y�z
^@�������i��%I��Ed���M�;Sj���IVb��s���%� \9(��O��is��nƋ6A
q����k�-�XR�<c�����M���9_N�o���U� �Ԁ�f���,�1�K�C�j���rN����^�X�f"�T.I�8�dm�˒�	�5s��o%
C�%��q��V�?��ْ�c�U+�8тq��3~~3�/����1y�Z�O����7���D�=�����%_&��1�/� �֫�<�qD��8bEvQ����I��>�?kA��k�Q$�m_���j�eEu�����
��%�Шe����WnZ�K��ff[2�-�^B�*~Yw�]�(�X��Z�l[�Cj��fdګ�bA�=4���Ʌl𧻓�h]*v����H����0���G5�F� *   ��_��F	�h�wZ�/MP����2�r�Ru���a����&/ {<��������Y�3���j���@{�n��S���0�-������=(�L�'
s��G�\!��!P ����:AMT`<W��;+]�1 uGQBbC���8Ne�l�o���@A�N@�T��Ӥ�XF1�n�%���D<��op?�/���KL�_"��qP$ųy����~>�բi7љ��\�����h����aT��	�Y��6�Ͱ/�?6Ѐ���F$�=`D��Z�#��a~@��2F̲N/��?YC�tG[7[,���Ϡ]��N����&��Q��k����QN�,u2�
��#LӪ#�p�m�m�U��JT></�+#u���ڲ��3��ׇ�q�7N�yy����)�.Q�ɻ�Es&{gA�Ū2��.�9	��*i�>_"L_�䲰��5���ѯ�CAЧ��̲����1ܬ��ʩ�Ҟ|N�+�l
��{�[��I��.L	��3D�Q�7ѷӗU3ֱ���uC�&4☏���Ut��:�:.�׺.�*"R���_-�-"XX�9\��6���g���ڑ箄���>7�*����d	!"�:@틔n�Bb5�Է��JT�X�Fρ��Aș����%��Ν{�CѕQ�ۼ���6M�ş����Cw�I��R��dQ�,����O�	��\��0֖�Gk�9��U�Jn8+��DB|Q�`�p�vDq~��f�ڲ/e/0�pU���i ��A,�[Y�����nm�v�~��L�]5�lc�biT������d�v�lz�.����nֱ�9;���jK��Ǻ��#S`��|�����cġ����Y�2�<��W(8_���0���9��I�Dʐ�%�SaK�6��3�!O�:�1�9��TA��w'�=�x����[ӲN�x�4�����Ȉ�x��1�����%K��ÚyFd���ԅ4�PB�T/<OU�Eaqe�	,౱�c�-��~�<U�ܡ[	��W>��%���TcWͲ7�{��t�I��ݮ=����:����� @��:��
X�I�w�&!�ir�ƿփ��p���o��M�4��`T�b��A�p�K��f_!]���ݜ�{���I��9�zo���q�Zf8�{W�a�x�sRN��F? �D���l���C
��r�[l�Y*[�1y ȇ6FW�Xe1(�mh���!�M6G(w8[>/��@{�xRo*���껄�Hv����Ah�t�9����X;[�K���U@�ޒ�W�u�S:4/�hM['G;��t$�=(.p�8��R��B�3;`�z�.aX�p1R&D��`q���n'� p�(2�K���]��@�� ��� NWXn�Ɋ�a.؂�s���.���t�&��O�"-T����{�Q~"k1���������N3r>�P.D����2�nB_������k�p���	�S�X``�c�� ���.�*XH��zI/�u?��&0QԊ��?�b�.9�H����J���t��8͌�G� S    �$�_��F	���RY{��4�p�j~����џ#�,}��Ii��8&T�v���xK,����C��_���Х��};�y����*0<G>��?�P�e�� LS���ת�dW��W�1�MD�h��Rk?8�č�L�-~任�*��G(���ީ�m���&WG���2IV`*$֔v?d�K���PH�܈��+��s��o��dj�J@�Oӛ����8�w�@)�*�	��;�	�?���E� ����Oï2)��'\4�E��Tϕ}���h"�O�:T��I8졶�d�9�@R��v����s��!+���QEm��	�G�i5��D?��)-��q �|�_�( �9�ͫ_����+D�UӇ�*�b儮�8o/H��Fc����1`�z�Z�`i�t ��A(�C�1�E�e�{ 2E�ȹ����C��`�"K���>��eX�8LeL� ckU�15v�����˘#6J������A�!��S��;��߲���vDZ��kz(�.3��s�m�Ϳ@^�c��!� 	[!��f9��I"}�27%�-�n|`j�W 8Xb�(#�$�s������	B��x��H�m�������W0��7Ͻwˣ��r�蔩��р(�8�����:U�[���]qPH��Db�T����8���7S��|���@kTͩ��>Č�� �3�$�/I�Q`|�J>.$�W��ni/�R���J|=.�ߗ�4������[�Cl��wpb�<��S����;��kQU�'���#���SC�:a$��w�L�����2H,�$h(����\Yfi2� B}���}���.CMs�˘D*��T��͚�9Lj���W��/��ѻL�w܇C�o��J�d:-tsG�Ϟ�L�/�����N"_AB��C�-����NCY DgW [/��މ\����]62�P�$�:z�%$Ӱ^Fz�H>�,�s14�Άe�Si�*wN�T�SXS���<c$f��bZ8��"��kJar�Ɂ��\�΃)�.�)G �t�Ѥ[_��1.�����*� ��=���29�"j�I���p���v9�rj�!�- �R�����P$
���0�B��Y	n	ϡ���9��Ȫ~�hB<�ҚSM�\jEOm�ys��{�E7Q�9/�$��B1{��-� �,�����V�.o]����{�cF�lb焢$���H�4}?<GV�L�Q�T�r?�م4pIXN�l�1�!n.Bk���I������T���7?�X�8�W����+[w�86�|O��%=��52��.�>X�b��<'�9+�բ4P|��'��0�l��6]���lC��[	-����9�ïۜ�gmMV�Qw3��}��ӹ&d��;�>\6����ޅ��ۮ;�Z��O�GO}���:V��s�w�Nֲ\,B��^��̞ﾊr]�FPIH��e,V+MY��>��lL�I���C}}T/�$��B��J���Hg�l��e�Ͽ�rL} 
�J�7
�1��|���95s�+����*�Ƞ� �	��kZ�۩���/`�{�A9zn�a���٘7�@o�Lz=��;�'Z���!