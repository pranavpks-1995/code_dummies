�W�>�\�"b�������*M �N�gWx���`��֕�s��NAm�V���4�Rs���o]}X��\�[3:ٴT��C}��ٯ����c����XU����*��O�+����-�s�)('�S��)�X��k�K�k#[�o&a�_�q���Dx����Y� %�8�	8��L���\z�;7���2���T� Z�r���׃\���}���l^�T�`n�n����9��tA-��;��=�L]����>'i�����ޯ�n���,է)�e=�w�<�b��1j�?U�����KȸXns,9 �n��
Ν�'�ug	��`L�
������
y��=�����_[�I=.�
?�a]@�{��d;c�oz���]o�Ґ5������ѹ
!�kX�$}�2o���֙
(��Y,��:t;��)WJ�LP�@M��d�'s�����@yLZ�}k����&���k��D`�*�RXS�+RtF�'p���;zB��č����]W�Buh<�@��W�!�d�7GE9QX1I=���j���خk����3:���J�#3iuJ��Z���:�c�kzf�y"h��ݘ�I���U�U�`[@F摥�;���s&�e�A;�EP[��ó���Z�XJ����m13�Ѿxsl9<$��XyH�w�eQ��Zst�y.E@�~���T��@����Kr���Tybu��sH:ȵ=� j�-0�������� �tET�Js/�YH���+����萀_�E$�"���f(X�=��������$ʏ��F���   � �-W���&8[u��6��� ��	�`L^�[}S�Oug���H�=��6x@��|�h�u�^<A���WLn/g�E����l>�P�?$�^�jZŸ!��ed{ոT�@�V�| ����m Y�D�ؙ#&�'�;��-	��!��TW�FQpG@�8{��)�b={���|�[+kmV���0��ٿ���Lg�v�\}�qiN�Z�����E�����7#�i07l壊
�c�OV��{*HgT��<�#��'��U�֋=_��$oO���u�_#7?���;��@?��v�<T����͍oxG��I�(�dH&�8� ;��F6[j� [�2�Q���*�;�d}��0��ç���X!�3�f�y	X���+ ����.����H���VF.�����>�(�-[F��tK���Zw���>���QZ���.�(q�l2tC� �>$��#���Xj���|.��)��nuhY���pȷU9��ś�`⭔XS��.��� ^Iaq�S�?��5l���H�;����yQ����țN�{��=2���A�)�d�b�:B@̟��2�|b����AF0��h�_��A}L�ɩ�p#��p٨�K�ZK��X�u&��b������(D�W�
� Ś4l��>yB/�`UqP�2�����{�j
�c�
Rq[M��b9�2�Z������~}�6���`��^�C�ch���.i��TM���$T~`:��m��V=��uw4