]�4��?����H�F��)�|��PZ�yت?��B����ur�e�^��g�@|j�����~-a�9&��2����6G<�}e��粧bQ��F�x<�/���%y|��#���*$�g�-���DBz�ZTC�µw�S*�jg���}[�9cyPa`�NK�>[a<M��Q*u����3���a(�B�&�ڻ�ě�F���S�o �8� 1�>^4d�0�R2�ܮ�GWd��j�޵e8ﻛ��c�b�u�?��$5)@6I���E��Rր	j!MM*��ZY5,B�1��q.?�oZ�Gg�l��c*��v��r��W͗��86�B���S��f�pl����j��NY�&4�ϨPU>�t�����Sd�eeFB�a�yu��'��B���   � ��-W��Ðd��r��o.��j~����c!������ v��%H�h� h/���Z�
�����w餅�� P���������m��/�����v�e�a>v2�-�C|8����n����6&=�sO�<>l����S2���b�ɉ����&�G�z�:�=�{ ���)��toW$���<� �m�	_Y�k�LD|�^2j�>�	Er�:���u�|4��V,�C���fNg���fv͂�f�h�YQ?�F�1��Ͳܠ��������{	A��Z��>S�<#����ՈS��kHT���gO�<N�AMO�8����5t�.�$�.���(:�ܫ���=��.�a��r�d�r
C�^�Sۋw{��B$��-V���x�/+�! ����t��J���5�I;R�( L�W�O�CmL݂Ă!x�_(��|U���r�z<L�����ؔ�^f�����Ty�8�n�	o.}����ޥ�����&�w2�=J>;���ɕ��ë^�w��(���SeҀ���6C�g>'>�W�����Zd/U���#��Rr}wh��gö�0&�ti���W�0���ޤY�.�bA&e1����_���ё��.�����g�_�!s������*Y��Q��}�6��`�]�����E����m�����ͼ`%�Zu��EB�&��������!��9�7*������r�<����e��U�� �3�,)#@�=�/��vu�O~�}�x��(�K�+6�dI�'�a�^����v� �)�aa�`1!������#�|�����l�������u/).^j�r�� tR`�
��HUS�-�NPa��j!��,��7)���%,t1��~<M� [���V1\+���Z�P��V�<�)������lɗf�t:xn7��[�S��[�+����u������p���������@/s;Q� ��
��@�9�����P��������ޛ{�� �> 6�
�pjj�2�� p!��-/Q�}�� ���\uk{?ߏY1_�[Ɔt{"-��}s��/$ӿ��&�$�U-~���~"]ʍ6
��e�I<KjZ*�Ĥ �8���! �
��Cq��d=�nzX�Jr����k�� {sH��L�7�inI.���q�������@  ` �� p!�� 01O�� �P�kN��%���P�zV	���}����b��"�aݐe��Ly����R�T��B2��Ϟ��D�}�%� �@��G��@��E L!,�)<;6�@��B�Q> !�k���0E�o�L~j�Y�l�;� d�0�0  �!��E�(B�v�@�(�Zc>m��Y{�S���h���K�g�de�k�!��c����~�ɥ]҅q������eB����{0p�����&7+s�V�P�����wy3��ڀ�H �`1B�R�A���Q�����E.;�A���N����x��M��Ff���Uʤi*��m   !��%M���mfX.� @ �u$�ʊ�'Q�fLE�����_D	���2����GB%i5��� �	J]��-�+|�2�B����Bv4s��]��vտ7go��������� ��@r=�
f�И����$��UTr��W��ٶ�'�i"��RH��� �!��&.�� XҀ��q�)xU��OhC�l^y���u�@V_퇁�P���|?�U� r(	OUq��Ӣ����-�{E3�s�|������ �@�0n�\H�8 1+�������4�?�~Y��ϧ�I3�L���)�.*�V8��VL	,��� !��%.fͅ �K KG,,|���5�����Xo��#�aIH�7��t�јM[�J�+{�1O��F@8�2��]w+e���}���ol҈�el��:g�| "���@{���"@Q�+�]*�