NT�cy@��n_�O��l�W����0YF)`���!0�ާa8���@�Gt�.���� <-UѾi7�ꀍj돭��Zk�woT�m�~�5���x����MQ�NH�x��t��h�|��������z����>��sHӜ���"r|�
���sE(0�ؕ�1m|a�Lׯ�����h�-Ėĭd�O-��9�(jGH++�E��)�◤�)��,nK��G���
7�ďut5��d���C���&���υP70*�[B�1A���@�bۍ�;\�mTg#�.�З�~���զ(ʋF�^B*��	� �d}�.�H]����Og/1�v�5C�u"�:��O� K�  �  K�*��]"q��|`��ۍ����YU�J����������Ot�t^rny�{�xfy��(%Mu��Q�SM�U`���;RLU���D�	%ȚFu�Z����o5Կ�s0)=��1���.��}�o=�IL���z�tޚ`~I̯K��uC	�6tP�x5�-s5��(wO>��c�K��D9�U+(m�o�v���7��qBC5��`\`�!�]����=��:�u��f��
C�<9�6��	���Ʋ����K엳p�j�-鬷���