Թw.���)��H�J�  �PC�x   ;�AK�c�jS�0L��1�*]�BC�,����wƇ�:ܛ�Uy��M�wJ�'�l2�:4dq��sG���h��E�S�-�w����i3�P�U�-��i00Ʃ�.���F�lV�J�tب�G� ۜ�|��LO�S�6Ғ��=a(���"�!�t�Z],0y o�bF�����׏&�4��C��n�ْ<(�D�X��f^�㼱B�o�~T�  0��F���3(�����rv(U>P��3y�u��-Uj�R�g0��D~��f(��D1����ъε��J�Y��z��p0���M�$h,���fn���u1;\���.���"{�Fj��P�8���>�w�Z=�!�`��8��;����?�1cmb�:[�
 6�1���
��S�I��-�G�#�@?�K����g@�v%�X�e �a/O*Ѣ;1BIt������GLZ�F2��};ǁ#�Ci��GSZ���i&w�¤�e$�<��W�Q�!��k�;�M"�����c�~r��h�0~���wqn�ԍ�זg޿�`;�fe�l=pӕ�Ǘ�T�{�?D���ΝA1ޢ��]-�/U�y��$� "�� ���`}���?�6%�e�R�����v{szǩ>?JZs�K���u�[���R��3Hs�"��N�A�����R�n�b\���P���l_�K �0�yѨb�c9#+b�/J!��b5v�T�����dQ��
�!c�5����{�������E��0<R%u\3S��AR��4���oҗnl�s�{��~*HY�S��<���T'3��t�J�A^�M2Dşb�x��6G�YZ�;Q+�bs�a�W	���k��D����熏:��H�T�<Ţ��
@鳪���}� �i*�`����o�	�L��`�A�]�lO������w'�z1ה Pg���X!	f�l�4mS62+�Gc%9��lG� c��:4�me	e��q�;��2����+P�*��4�}���f�=���H�<E�/��e��J��!P�������*`�{�MU��I:2Ǧ�����1Z�����V�bfuI�w�T|kV�����f���7����f�o^P�p��h4)Mb�,��ed�5�èaT�S��-p��y�G�
�1̅8��U$�!#A���bB�9��0άY�2"m�>���;�Ыq� �)�w�$�>b�6�i�`���D>�vDђ�K���%��}@����%!:��34 Xt�\���6�NTϻ�V�q��I2�jB/Á#��%�T��y�<����`h���{����¹�GސM�nEu��q�L���T2��Gy�ſˤ�?�en$���t}HT�x՟���B�9U��I^ʪ=�x���e>5.��o̤�Rq{b㰔
�h&�����dËn�κ,)Eg�L$k-�!B�F(�e����^@����j"DNK��0�dJ"�B����u�?�~���닲A��0�	n�!,,��h!�$���x���ߌM�n�N�����3fR(��8.�P��,R�<Q��ê�9j��l '�xO�G	����[��<I/L�z���n�}�t�z&"@����r|��.��!�S,J_	2�^T�����7�j����$C*�CQQ���ߎn�[W���Q")��K�+P#��\�M�c���`[�2�9�Ll��BP���D�	*5�nI��p.zS?r���{�.:����8Bg���i)0L~��)Xu�lÀȍ��<��Cd`�t
����$�P�8��E�;	��N)pAg��J�`B��(�?��7W.��v��kòR�L�]/��@��:���zӕ)�l_u��>���8j���D��o���T��H�(ǎ����5v�X�6�6,�ni_��_$�D��P"1��mf+���#�K��^]X��a>�d@�X���~̀�O�QA���/�¿kD�ЙbRcC^/�|.�(.����0y댑����a�{�M�	�H���5�1�1LL�̑�_Z��X���Vg�cN���\��{�����Y�7/�m&S�;J̧-��]���'���o1��N�������#�Kq���(}+0f�k;d=�|�-����3i�溚��;�9d�%��}�P��#��\� B��2�,�/�l{6���v�13�	�y�%$w,��@௥l]E)�	�(6�1h�g�q�>Ύ�\H�cqT��k��z5��͔i�i/5�Ԍmጼ�&>kN%��A�$��W���QA����/gh�2��%��LBZ��
/�Z�MdfeC}�Ҭ=���VZI ����5�=%����5%�ȃ�O	�L���e*�I��&�W�y�E�?6�cd�@h#0S"R��ytP��k�ug�����T�b�R!���U��]d/�ԛ3�h���l��g)�x�>>{��%����R�w�ƺ"�~ۿ�.��e���Lܖ�N�P���(f�)�E��u1w�ٰ5�������d�;p�n�;l��F!�8c���+�Wl��R;��:��ˠC��֨}�S�*v�{j�Z�q7���v���Us�qhC/�y�f��w�r�	Vذe��-���S�A��=���!�	��4x��֏e��\i3��� �]��&i�&�2$�w��4�s6����҉brP�~�iK�V�aE���I�Q�ͤ)Y��	�FB稰����x$r�7�&� �T@�ti�M�-��Ah�vQ����r �t����ӭ.�#/�F:K���W�U����dY&M%?G�n� ���w���Xw�\���kG���>�E��q�B�ò�n�"U6W�y�'Ҏ�(�@ �EO�&�ud�x��b���2�/u��X�]���a���#L_�#���x�鼑��1���i6j�j�2�9G�����>@��2m��� �vM ��7���ϮC�7*2l����Tծ��0��-��?˃��YD�O�I���. yf�t�J��Oz�Ĺtby]G�Iu��9��m�thf��ݚ����TT=}��p��)u���7��?dFH��F�i��˙�?i����pذRܿ�&Ӄ*gT?�$�^еP�9S�~I�q�~,6iOF�6!]g��)IMy=�܍�ϴ����� �Sb���j)���ĒF]���:BM�֕����.�q�l�������G�{bx'zX�=�%��zeںa'n����BU��9���w_nrW����Es����V^�>�$�d^�寋�����q押�z��F5���inh�mySF�J�{���!@���T��U�;z���"빸i�]���H3 pZJ��%(u�"Ԑ#8As�΄���p�H��T�'�d>���xĭ�o�R��V�����x2��qP;u��W?</T�;�ҳny�����A�E�n���η��}������ԿφR�~R t6/��שݴ.�ͪ��u0GC!.��+խx�p�/P+�пv_�bS�X����C}f�_���I*S������VL���; ~さ|��_�@��&Ȁ��q5rPg����K��"=��v����#b8c�/�����ޜz�/_?k&�@��PL_Z���6��_^��^��"g�Y���ї�`P��͡�����F.L�f�-����2��@(�~������L���{�ځ9��eK����K�CvD�K�=�N�ɻ�l�S�oÙ2�ei?��mT��G���[Y04�Z��"J���:�J$����Myi��}���&�K�<Ii�'�m)G�9�������r{)/Q:$5�����L�����o؞�����6�U�9
�i��5Ҭ8��|P*0�]�a+�`��B���|n���K�wU�~�o�q�f�o�U�Q��ǎA�H�w��;��a��	�m~/���|�!���k��ɇݘm>ۚ�P>H7f<����^vXd �5e�����:�|�Kؘ��>�Z�o�s�J2���X����u���Ĵ��i��'�51�8]��1Hd '��&�g�c#��� ����F ��Z����I,����#q��\�AD&Ԟ�а�����JO�~�q��0�|Ng��s�K7�C�a9Я~���E�$  ��ĝxc� ��K]V@<>@S�BX#,W�z*��~�4'7,�\��ƴ�j�t~�{foD _!�e8�.8	��z�͛�
ZҙH��15����"$|�P��jy���誹3�m]��',��+"�^�}' ?�8�dST�����]�V����J�+��`����W(��*�w)'vC�X�3S�^�kI�ܬ���Ҏ�>�-s�!O���L��F;A�v�o�����}���u}�;�6v+*�>����n�WӼ����l8ν*���Z5�����V�-���Ǒ�s�;�5gP���ǜک���<����f�el���]r����?$+]|�AO���@������w;�<.5༑4�� 𙫵U��tS������	/�֖���M�A�Z"�-z�<�<�+����g�$�CT��&���"!>�h��c�WG,"���!@9c�d�xvnƼ[��6y� Q��t�q���T<��״{b�5?�������ο�{��sW�t���+�= �a���$�C$����OV>\�F.%��X6z1�(����R�PWF�X�?���${�f��A��,w(ct���A���O�YNz 4̉�׾г����O�(ǲ���@�V��"�	��D?�ɢ.��_�.���ŌF�/�������q: ���6�<�oB�g���rcL܍��zPӃe؄��e\d�������)|UN	����&8ٷ�)�
�~7<7�,_���?�I���;�����,ّ7��(zݪ��3�=D\��D�1�3��L1G��
;�ďޯ���{��*���IK���1�yb_���{Y_Z�m.0n���Pʎn��j-��'�G����Jq�j����ah�=?��qcֈ�F^�1#����Ʀ��4�ʃ����	p���h>y-�~�2Ȑ����mq2i ~Q	 zT�<��g�p���������*OOa�������*}ܑ�vh�+Y>�+��W6Y����ӣ��Sq]aeo�N�k��;�EV�R�5J�N��A�	xuCXa��"e��":������-z�C���v�F��T����W^x9��S��)YnZ�=,���[����].�!��(؀iPw`Fb�=L�v{m���I�=n���9�~���B� C����6׷ߒ���3o�'����6�w�O=^+�>�K��j��;�s��%B!Bn���E�V� 9��k�Ր�.I��&��5<����WJi" �Vʀ�����JB`�Ոi��}9��L�[��9�YQ	Ӹ���D_� �  W ���_��F4B&Hi��`_��Q��j@Y!�����dG��˝�`���e�§E�Ը�j�6
�Ŵ9L"�i���G�a����u��&u8��]ixZ����V�
�ĭ��n�R��Hk\��2��0�!��y�y��)U�J�8_n��`"	ZE����%ǩn�����ք�����!M�JN�tž&�	�@4)f�@��B;�T�/�������]�a?����ܳ��EP���^���ڛW�����j�=<�n;����r��g���p����%�t�u�r	}�ʢI������j"#�:��ۚ����Y��$E��j���(y��b�������m��'��C���<jM��̆1Q֧EI�bh�Ng((KF��d!_V+��~��&��"M�u�	�3�,�5�y��ݸ�"A2M#u����l6�jD_�"� �쩩!���E�w�D���!`�_m�03��+�4�FB?ۛ�4�����6A�@�1�/va|[V�s���w���:������<8�D��O�^�����(֑��jfLGU�`��`�$l:B��a��Q���h��=y�=�z�ছC��*�{�S�n�>���A� ��'	#�-���T ��}�"�#	Jil�E���`3T��2�j��I.Dv� ��$<��#�Ž��o�Z:Mr<d�͎�3���G�ax�BK�)SXmHP���C�:��h�I�N�u��b\�5M�ZL��ٍfnC�2X�I,���Z��Vl��ݲp��!J�%����	�݅�+%�+�5������n��b���(̽�D��h{a��`�����	S�h@�D�㮅��n^�4��M�㠼H�AD�k[k�(4 b�]{۔��a)��Ӷ����J�-�w�@u�B�S	~�7��o�ؿȧH��x�&��t�=XYd��C��:����HΝ��ϯ��hD�PԻ��m�U��ъ}֞�tņ	��u ��%H�pэ�Y���$��rMC?Z�z��g'�B��]�J\΋\4=����A{ o���BFvH�c�o����v����w��V�]\�L� ��=�-a�����g,]	�!t����Cҁ �   � ��_��F1N2Hp��]AF�Rfj����:�% ��)R=�(!B?e �9o�C�4�>!]��(�LpMܥ}��������0%V�4:���݌B���#���卓�@n6�Z�M�c�Gq��,[�hNi&��+�ȅ�E�����^ǯ��`K �}*`MU ��jL���װHLh�P����E��������Z{�������\^k�(���ZWd~�f}���l/ЉK~z)T�U��#� �M��R;]|�I��,[LN��$�^;��ׁ�c���u�o����Հi�5��cՆ ���@Wl�P���c���9�=ސ@���к�_F�����P�jb��-Cz.���b�"��$��X�W�.$ID��W?�0�ɳ�09W:͎�����3IL4�F�UX���~��ji^HE�k@m��FJ^RI�޽���:o���w�J�N��j ��Ɍ�Rݠ�������2�T��[dPE��k·�
��Od���|N0��F�)�2�� '���{hG4�(�C�-�'D6��g�²��O(JUEx$5�M��/_�*-�$�R�����y�ʠ�Z{-[�,϶|�D��QϮ�DQ-�J�R6��eQ���ʢ��M�5"�H[��w%�����h~���m����V�ԽD礪d�(�g��B��)Ơȍ�׎6�T��
��qu���|�2z$�-���tz��[){��/��R��;Ǉ�? ����S��G�4�� 6��'�J��Ư�b\���zP���K�Rff��i=���fҒ
V���ﬤr�j���;5v�?�{�� �	C8�}� rx,��P���I`��TL���u�״x}�M�ь6
o@�u�U���̿:S`��;l�"���~EsB߂3�{�h�Ӏ�C�]�Ҽ� �t�5B�?���3��ת�,�NvNb�$�B��)e�/v�o�Pn�~�����;,�BŁN   � ���F:0枬Rv�)�`����ì�B��z%�Q+!_8k�4���P\߀���'������Tn�1p'����k�d����_	��d3�"x�*e8ʦ�� ���>xQ��w�
G��,r=D��~�;��'�8',�{�ڿ���
}a*r\V�MZ:�p,|ٟW�Z�`(�@dbBuN�^7�vU0Ҝ�(�{턐[�}����̏�����E��\�I���Oz�҃"q�ɑN�y��t��n�l=c�� ��bl�+�"��1{ݿ#���lq��X�D��f�b�Me5����ǀE+ĭ��H�X���<��):mQ{�jE���8{Z��)�=}������U|&� ���)��V�[Qm�z�,Ѷ�z��?L�[,��@�$��YA�uʂ�	-^t����1�֎w���b��	P0Ko�8��L~��M�����Ϲѝ#�C�G[���n#��`a��:�kv���
H'�z���d¡����]4e��0s���6@y`��=u�t�B-�O�ʔ>�{�ʣ�ם�H�#;xJ��1�eOŵ_ԮT9(�ɏ!0�ƈ�̵���>��F�'�}<o�fj�_�Q���Ym݌���ʮ�U7������4Ҏ��*Թ
��W�Ҳ�M�xi)����ΰtp�Y�Y��WByڒ�55U��0DF6���O���CZ�k܅�4{u0�!���K��   ��P�W��c���OF��z�@WL������\97�n������"�Y	0sMEg;M�
�G�����.���w��]d��Ƃ��\Ev���dBA�\<�5��i=�����bӪe�)(�5-@��W
L<�N �G��m��\�����e������*^���r������G����OϹS�<|j�u]�Ġ~�H���JC�WN�J(���4aTk���t>�����+��"<j&��ZP,�5{?�H��p�tiF�+Ў�)	�`�X�\�R�N�Y��Y�������(�ߺ���G�X����T�60��S���a<M0�"|����S�H�g'D7��,ܦp����t����8�9�o�ǋ�c������Ki8;
oY�J�lʛ������7b�ie?�*hF~��<jkPơ:,bs:�WuT����|E�i�p�_��;KX-�'��D�un6�<l��2lr�.X~8.�=���y��H��K��o�?���X/�8S�m`�괂�����x�Y޸��W����{y[��f�^�.8��R�����#���!�n�0�okM���Uw�� ���b��IF����ot�n���<��^\n�����ƫz���KG0�N����^lM������9��B��uyz-[���tc�R��,��z�A��Ȍgj�6���6�:��n)_p�IV�_�ܰѷ�ZǅU�9�H�7T��$����\*��+\zP��MC)hTfX�\��V�O�䙰���ɻGW�Vꞓ���M�P�
G~{�;�<~W