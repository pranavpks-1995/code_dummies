��C��-��Zd	̯8�`兩k|�Pߍ�H��\Wτ���
.D�v�-��y2�Ђ4�ʠs��➆��x���f=�͗]����<"v38�4��|�&�}.�"$�g��k��ӥ�ɖ�P��; �)�:�r6�_6�v7�a^�q���n�J����"��3�e		�;Ζ[�!�8%K=��c-%y�έj��z`�@_y6A�� 2�x_{��P�����:���Ը��D�xw��$�'����z[T��+�1&�Si�'��ݦ��*ʩ�s�Z|��@��=�
$��`-�`�6_��ce�R8�IT1���;�c���<`�k�x����y�wH)�أ�%&b{c|?�����j�!\ܑ�p��비Z�l�xo&�4��»��h�+��N������BY�x��o�u8~-��(��]�o4�J��<}�xAj&���F��W�MX�0�N��c=��n���֑B[,��w��+mv�~�zd,���6�?�BSR��k_��ӧ��~�0{�*�[��*���JPQbz�����d�'���%�R����F�z�O���k��"��?4-
�R-ď%�\Ž7���Wb�%K�:�!L��`�z�0]4�+��n<�z/�+[��-1��Ο
�@�i��6c���bߣ�Ρ;H=��`j1�89�����m�������0�j���C�G������>�k8IlO�֡��VCU����ɯ�|�'�G����,��K�k�WOm�cW��&��qb�}Q�e{�}.vw������� �!�\x���ߵ�hs��Xv�T�J�Y9���tC�x�g�
��O+ ^[ekuT��R~��&� � �7+%?�s�&�P���_���V�mr�+O7Pr<�g�P�U�����^�3��&WF+X5�*�Ǵ��o��I+8��;R��s:��"��E?��%L<�m��.�Ow\e�cWt��%��a��r��l���=T�4:�Z?s��0�+E@�i� $�H��,~�T]��ݖ�	s�;� L��
q�5,�ɩvǬ�ΏSH�"��<,q� �!~���-w:lѣ�ȿ��P])��hx��?ۛ��*6k�q&�C�Vw���x�����`7��yfr�`��%��Y4�S��3f����BbJc)�͆CA�t���A�`�&4���޲yl�%�鲒��S�aL,��W�[���H���Xm���z��~�Gz@�/^�x��1"���8�C�}~r�Ȇ�Ky>^�2M����A��\����;�ߓ`QB/����aY���r��~��`("���aYg�~���g��I�Q�1��L6b<����Tk��H0�qn�|^�\��*��0� ~�_�� ���	�N��~ 2��`�X-匒f�A�7Ћv�@����˭��`�|9����"��.��b��Kx��Bh��!���k(�F���=}p��K������a�-3�6�&��k���V�����^x���[��'�L���5�A�T8��T@�'8�ϚL��d��/�.I_�x��k������lbP:\�����|���qW�hĔٮ��r�?
��Az��Q3R�o�Kp����W���s�IԦZF�B�ۀ�� e����t~Y��ןT�G;�4�"54v���
�{r�8��Uy`���#��B9'�C|�p;.L���jY�6�	@��ؗ���B�ƹvA5�#��I��ԥ
hK�Vi8�c���+��-f`�sS@�a�
�V���C<���|�r���\���)���X�_�S.{�ލ�z=��.����9O��p�5��r�N��<#� �랂^��1|�0b2�������҆�uL�H�=���P84|�[����!��Dĩ�V�Ts�5�W>N��gM8@��rd9����y\8Ȃ,�-*�/�bGM��qx�w���1ćj���φ�"�6;�
��ְ*�$�Q�,5�A���-��p$8�yC��E0Ď����$'�f��%�f��(�jz����G.l��Y�� �����d��I5�v6Ev����~�� �@�~%Sr}mq��������	zk@Q�Z�x�s�}��1J����@}:�R8f+!�r��-�1B�8'wg/X�����y��iH�~?�J�YUa��P�l�f4|JYs��ӻ���Ɖ��OM���/�Ck��t]���*C��v<�y����>�E���>�%{�tb�2��}�M��E�)<������o� jQ�޼�m�I���1~n�V�3�prE�M&yE�������Z��ń�D�OP�t�S7VJ��)>-�6pdx��9!�ch���m�A&�#6�7Z5�m�+&��w0�2܄��E)��T��З`	����〩���L�;!�L3k�y��e�es?�lD`"m|��LP^#�`lwW{�׫���j�{bP����(D_sw����u�r̀��N��?h� �Pm7�NJ���������HP�.�P%�$]v���ʌgk���$q�4W���/i��&�>Z�k��PW|<���1��*���`�P������IGGÿ�/���Bi��  a��'R��c��Y��o?>x�xŨ�����i>,t���������V��!�@Q���2~t��d���+��2�q�AL�x����%`�d��h�f]�*M��I�Z�����|��m>T�}�c~�:��H'�'���><�^b�2�yg����E�*�D���1;R
ó`P�Ӭ��=	��
s�ϊ���S�S(���Dɏ<����1�V3�X|�O�~f��/ĩ0쵮�p�UgW;����1Q���.�^������j�^"�H���W~�g�s���Ԫ;;O����&���r�,
��~Ӛ�ۻ�̜�$8�VW����
�<�����î�5��� ��\��Re���Ժ}��	�{�:�]�@����$ǰyˏA�Y����sTU�[�>ñ��|�S��ܲQ�L���+�m�E#�jre��1�g�aYpK�~�:��8v��ۜ@u:�J���j��aW"���u�O�0��������'���:_�����KZ�Y�
C��K-�(bKFq�]��0c�Mp��.Kl�A�2U��0oH@g1�d�?N{Hh�����nu�OӨK=�]$�b?,E��Ϟ��A��  � �F�U�z	iJ�F����'� ��� �GnU��]�M����E�bS:#$M�
�Ϋ���qL����:��?G%��{�BP��l���,�+�;��Y��ث�C��6�>�V#ܡIo���m?_����nK]W
�n~UaWY�0o���|l`��N�$sƶD[.{�.)-=�(��F��8z0�K�~|�E^;��G�sE'Ѽ|�"$]I)5��Y��D��m��N�H�X��~,c�Iݎc���ƶ�0���~^��r�MDIQ�X)3�����.X7KU��Xލ�b�(թ@�0jұ[^�:P�o"�DPߵ@gjI؏z�+|�(�}{�k��;:�'	OS��	5��Y'��De\��G�<�e�$m��w8{ޖқb��J&\.�D��۶ ~@F��&�A�zW)��� �AX�ـ���t��#�WC��6O�e�R�������� �HZ�#{���L�9��A���   � �f�u�|*G�^�Y��@k�O'@`y�/��P�o,k��� �~��\�=��m�N�m��'ͼE 5�e��@=�;N''>��Q޳R|�|���˒x�9&�����bT��d�Qf˪��(�͚��0ρ�	����'?7s���,g�}4���J�5f�<_�d�gR� åC #	�"V�BZP��;mI^����A��;Ok��'�L������&>�����S��|�@@q�k)N�fmBh���r�*�hʶ�S����Y�Vos�����ng5���%� �Y#$��¤
؀.�K�5�$�ٛ���1�P˃V��,$�Z2��d�OU��[�^R�0���!	�B����>�n�#�a칰 {�r�a�M��Sg���O�?��U�*��į�3G�r"#l���` ��\ې��P"�3���A��   � ��-�����V(�vI�&:�7�=�m+���>�k�F;d��\�?�Wț	�F�p�co=�*+| ¼4��W����jq��z��VW��l�^ɰ"F��m$����l�ۯ?݈Z��4�Kx�k�e��WQ�XJ�J� �!�)�q�0����ր9w��^]��o)�y!e��V�o�	��+b,�JHR�Q�<�C�bS���&�g�?%@}:@�!݃�:鈱'�Ӵ�.'���/�܂$� ��>{Bb��O/�I9E�'@{zo��jId����uL��g�B�����ۓ%����՚л�լ���h���5�C�Y2�1�c#P�^4��a�㴛.E1�`������Bnj���I'�b�0�&/a�0�	���w\��K{�8��D�X�x=�RN���p&�AH�VL��   D�вU��D:0R�!C�T�	G3,\��p�Do�5TNy�n�P<��3���Q$��N��ⷿ����a��Թ>��e�����s/ $iR�I2��X�!�%�+FI�6�X幱5�I��c�L/��Z''4}����Qy3 R�P�D�I! �F�XH)�Lv<�/b3��?J��w�`[e�ؽ�mS��y�\��J�dÇvl�P)��̈́�;\��5��Z\��V� 3Q��V�����Gԙ�o%�H�/j��c�a0b���Nl���a�8���7}���l�L��#�̖��}Gx(�(�4��l30\J�P"��feo�ד�ץ^��d<1�Eð��D������8#p��9�yd�&̎�����w��$��W��B���5uR��r>�e*��I0��sY�9e�1�f�9\b�Y �\��*��¼���Gi� �w�ȟG��Y���KkcF�W�.�����0+�Ƒtl���rL�7zg����O1�`,ȏ��\�^or������n�ULag�΀t�;C�R ���%�~�%�`S��v��y��!\��<�1)�w@m�.!�B
��vN/�C$�	@9� ecz�4�� �h�"��rdH��-f�(�d*,_n��&b-Z����,�zİ������L��
kc˵���XBnI����7�Y�0\�;)8J��&ul�������v)�٪�N]�~�i����W�.hZ�`��Ӵs�k٤w�����Ս�g7���І] G��)\P-�����4ϣ��=��Z�?L�%�1Pcg�,C��2�!���l�YF�'��XT���fLlm�H �G��[��Y�tk�j��"��5��&�:�}��ED����+d��U�q'�!�h�\���	�R&�(+!�щ�0G~�{_�O�8˰%F��#M�?*���xu�;����R������I����㘿>ފVL�G#(_�M)[X�D�qV�<��C��,���ӥ�G�7���>��HK|#�D]0���2����Rg�xI �扒~�������U�k�KN�Q���S#�R���f���S�Z��ǝQ�ܱ�f� +�3��*�^3��P�L:C��P/�.&��A�L~�����,�悘|u�1���eq��z��"�޲&���x0T(�@7+�(I�*}���&�nD�\���,L풀�,��u�GL��۫�2(&��[2"��wN�xm�Ɓ�	ЄB|�UY:ǀ�D�
Q���4�����{�e��#v��Y�.E��n��s��:���u(EfNB���u��H�h}�[��v!,1�=P �FO�\�}����ڱ?��on7���\S�}䜑�Y�miq� ,�c�3�3b쉩ȸl{܁��<��2Ε��ŷ�oc��/Jh�j��5���x�3�+�|I�*-X�-�b3)�+T-q��E�����x�@�Vy�����E�=�>gn��"J�w]�p����z�c�^�&!5��I��+�;�sS��`�^�bR�ͅ��f{,=���э�������$����Y- ���YY�R�X�/ǑОQ�c匪x�)��>`7l6?�8b�F��&)S��qXb����IcRI�
!_̭F�N�x�9�$y@#��zA礢C+�}�����S�[���a�c[X�=EjH�x�(��`t���TTYQfۂz-"z�����6��v�����#��Vb�xxF͓xQR�J+�n�15[Vn��i�g�DǵG����mėǗm��?��Rh(�4fy�!�ӻ���*%��9y�9.A�����ڸ��*����R�_�
N��G+�jk����a�&px�٠a�BQS��������Ͽ��rhR��(q,�Y���^wp�{���O�/ko�Y+s�)��!C�~���ZD
�����Nߓ�g��Lv��Y�4Z_�̰p�3��Z��:>?�B��Ɲ��9xTҬ������t������$ʱ*��2C�9��t�K3΢&�V��Y�����j&d�S.r
�+p��G��5�%�E������D��
9�L4�4C�Ls�Y��e�'z�n�R��J5��'>~tXwU�h5����>a~��.R��'�zW/fw5� �#�-1=���M�r
�8���L2����H{	G�r6ࢥH��?�w~�=B�Ä����D�;)W>�mUyEa�o�Pƿ��ђ����ՍDŞ�(�
��=�F�Ws=lc_��.r/ |E����	�JNf,H�wyaB6�g;��sN�L��##��̤-2}�����0d,����fWzv�� 9n�ul�C��ZiV������hɼF��=��W7o5��]�"�J�o=�J�)V_ֵ�j�1�t���Xiض�[�673CS����4�??���i<�'+�O��?#e��)z��6'�5���(�)LX�I��j��갈ź����n����/7>>�
F�{�Y�7/����-&m����,$��&�[jƍ��]�LnA}�H��jF3�
�[@>�ud�;A��Ϛb��Ѕ���Ǜ��Y"�@P�5J�w��|"Ƞ`8xF�8�Ȕ��{-LZ�b�V�U{�A�W�"�z��������Tuk"�ƄS��G�Ve�PtCn�0���*d����fN��"��}ܧ֥�21h�{��f\��
զ��Y�]���
��:J��y�?]8�<FZ��U�f����\n �<��ܜJ� 7�W�ஸ_���`���n�ș��Ek��Kđ8q�(��\��c�~k�@;`^۰��bs��Z"V���Aj�z�Dξ�#��_�A���i�x7�=	D�0n&�E�'��t�G�hē��)�v�9h��JN�̴�f�f(�>!���u9�qmpd�?�����L7�Ӛ��fLl�n�~��ؾ�\����?�M��U
��5�;ʯ�>�T�G��89��
b/��$���4�T01I}����1	䢽�X[e.o��J2�=%Tx''��Gu��ث�퐞�W���Z�;^Zz���� C�0.RU�[�@���6�4�!Mx��M!�a	`.�i�f�ac�H���1�8�Ԟ�J{bU��:B�=`�Z�?F��������c  
��[BA���g"3��l}��"�H���2&�W���dD�)�hz�g@o2��w)۝$��3��x�G4r��{y<. ���7�K�G�H�
�k��ă �}����&���ŏqB��ڦ-�s!A.�,1��@6,1�w�?K�K<�_L�*�`�����#��۶t�;�[��D��p�J>����Ѽd�K2d�{���Y'��@-�-����<��e%_n4M4>�˿e�L���d�э��Ҧ|��=^a�kQo���<����&�3��#Ƙ�*ΡP�@��g�V��X��Y�x4)VqD#�1�c���"���K{���/FؕE����Jq�ڝL����]I��p���\�g'���>!����É(�,yŇ�tH�<��c���O�?���v0�7��JE}���vb��D?���|c"����&����Qx9�#l˘��M����>��#�T4LJ���� ��h�ϋ \  c����0��R�e�B�[�Gm��a}~����Ք�o.Z�x{�+�-�R�@��1n�~���d�o,��x�I�ST��Ӳ��^/���g>�}�_`��xke$�th�D|ǧHke;̥�������0ekb }�2�fM���4]���\�-�["���ߑG�z��q�����`%_m����c?U��R��*�\qE.Ej�T�#�����ʮ-�� ��8%?�]�~���X�ĝ}S��q�;���)��ǲ�s�nq�B%�S�K�C�95���pʦ��\�b�EP�]��76%H ̪�J�fi����}lg�/��$�}��;�\2�33�1}�2�n��O�V������o�,T��_C�Z��~���7�\>ʟ}�l;W�A���U!�H�ߒm�yJ���R�[c�E� `��<l��%�ĕPZQOT���#�7��1>���s�X� ��7R#�����%��U>*��o�E����c�sw��4S��c��J�]�������?rW�I�d/E��a���͡�k�>UZC֖Gd�R�����&S�m<��a+��e���:�8�N���O��\O�G_��Ns����FIӖ�<����:Kt}�X+�Ԟ;fޒ(!�<��)~=�8i�	�nc����'G�ݨ�ST�쯓+2$��o뇲���Y,�|W^+����Gv�?;�D��޶?�G���VC���|�~�A���3�fאa���j~�T앚{��>��7l(��(��q��%#����gD^�Y���}�p~ֻa��}qd}4�{�i�̔lo/��{]:'�̰YȖ�N�w��v�+�J�~��i