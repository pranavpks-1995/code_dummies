���Z���*.v_�xG��$ёjO����Hx�J�g=^B\]��y�g�4r 3E�Q6|�Nvq��ӊl|E���S������/���&�7�b:M�n@����塽Ai��f�4����R�����ơ�|���ER��؊������W7ە�	����qLb���_�"���X��w
��'���;�?)O��E\�q�_4t�y�K��t�?SA�C��u+~�`kܭ1N#�?��/AyY2�U��,pB[��V�Ǖp�$�6W���I^�<�f�ⰹ+E�=�*�,����z�U`G�h�ACy
�:�n��z�Ļ��8�	eZ+�mV��1\�=��|b9s�^�_�js���l��p}dB�F�AQ�W!��xh�[�i�Bɇ&JE5 ���gv{'����ɜ!��r2�#$%a�I��$ɾ�.�s�Lp~��I�}�%!5�0|ap��������)E��C��rD"Kf�s�xB�\��;`��@Ɓ��=+��:;=?l�-*4�j���	@��?}\��faV��@�W��LC��w;�.���\�Q���y|�=���\� ��,a�@�z};0mI��=FY��1}ɡ��r*4�N$����}��ߡ/Sp��m5�0��ځ��ѡ���eQ>�叻C�H��Q*T��_��ǹ��N����w������s<Z���4��c/,ޘ��)%�Fw��������t Q '��]�0ݜ8����jh�L�Ԗꁑ tW(���p6_������\DEU��ۂ�	S�h�}��L<s��p�qI�CɆ:��^�ep^i� T4Csʿ���N��r��r+��|�#	A1���8���(��c.>���%Ӎ��U��W33�	_ОY�Z�am��Vc#J����,>u52�K#�)�$z��h����6E�&?�,�;���H���'P mF�R&E��4t��ڣ�#