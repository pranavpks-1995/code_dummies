�6`���BZ�
0�ǃ)����A=pA�/�\�yR���1�Zf�4ێk�W�M"bJ4KG%�6a���k�*��C�Г����dp║o�$ర���dn�"Jf5��w�e�k���Ș���5E�#�ۣg��Ӗ�v�:�ֹ8��ږn� 6��Ѿ�n3�o8��~���~C�朣�����_Q���jZ�k�*T;C�1�B�d*H���p�'�$PH�t�Scz|;��
W�>abq����-��.i�QNՕ��?�!kʝ�w��6C�����gݪ�-��ىtb�T|;(��-�^L���U\�=\g&���f|eYƉ�k��0^X��>��0��K�mf������ϳ�Rp'��A6�3��>�pݽ�c:��؝$��{����N�{�tU�DY�e'n\m�έ�̄,2�kLǛ�������a�7�b3�7qjX�^��z�X�I˞����]l���3���l��;$��=a|P*���,@��mz{`��=,��̰d�OXx�>:�)g���܏�l)�u�5�6���%jl^Rvk5�3l��Q`]��; �[Q����K�q	���QY\Ha�ª�Z��gA�?�l�3å[��:8��(�Ld	�����=߈�w����W�E3���I����ne�@���4H�-�WM:>I�:�Vm�n.��O��ķ���X��r!���M9�7y૳_:��ܙ�錳©j��W/�+[��}BuXu�7L�|h�8Qs% �������9�oCױ-���*H[�~�T���=P|uz׭�qY#�E�P��R��2�
?�6Xl�CP`�h�k�0�C�wuIj@B`IV�_�A�m��P[}���2ŗR։�n�kB���d����JM�6XǬ"��T�����g��I�S�c��U�$L��6���%'nLc��vo��t���Y�:w�x�?�����[9� �Z��#-�CB�A���xi��/��l�q_�4�qF��ę�r~��&@%�T��������tF3�,�ɍ��;�6��Y��%���TQ�)ш�u���z��@��Gߴ��MN�9='U�~�)4;�#��@v~�����g �ľB��ʔ�Ȑ���Q�k[1]�9P�5!oMŻ����eX(~3���q&\��6��aydzS�5�(B��ܳI>;�9k];�S>�<,6��rx#Ao$����q�qA�a�*j�䝼���;�V�u.$��#����V�Z�V_��vd�-.��"Bhկ��Lw
�p�%��j�/�pIbrz�&�8�P���`�j{�>���OSy
j�.��j�~���9<5�$S�">�he�\W�B��c&ޜ9�#��т��Na�cZ��+h�e< <�+|��9�yV����t(>G��&��PV��Ew��#��b��Aٟ48)d��i��.K��H�:Q�I���}�:��m�I������v}�5�n1��
Co)�X�:s�z�I�8�`l�Q��*:Q$�l.�.���2nѻi��f����}{���I�i��w�ݶB͸�J�Y�4(X�N}A�ku��S�(��Q>R��V犚��:P
�d'e)�F��	J\�w���J�o��!��cB	���h�Q.��f���N�
6U��#i���:H��A���