���v\����
�E�������+Ș_�a�"����� 5��I\���� ��~���<KT8<N$�V[p�e%�#��zs����\f��S�Q�X>�2#��2ԭ<"D���M��sG�;�$���������mo�(c�:�v:eOEvP�)�������"��H)-�: �;��qվ)F��(3O
`��7|4��ٔ?ӷW$櫲p~� Y��R��ljQU��A�x�>*��վt��K�8f�mg��Q��$�w�X��Yd�$}�X�5;d/k���﮽I�sc}�P�1�?�A�bb]p���!t�JZT����Nj��T#��ݽåO���:'A����j2�>��1	�G��;��R[P�H�lA��4��4|HD���]��}��b��~_KGnܿk�<?�MY�.��l�S����uL�!�.�� �W�@���c��"Xߝ; ��������(E�	��$�@!c
�.��
����S�o8��*��Oe?!����5�^�T"�?1��NIsi��FOd'I�)��������#�-�uet�ڋt��8w����OJv�6yJ>�j�N��e��p|��X�������d Z�c�Cp�@"��aqr�=M�F�M
a�,�f3������Z���3��Sg��e��i�K�^�K 9	�ѯ��"�v�kΉ��tB������#�X`����R�
F!n^M�§ԅOY�?�L�L+H��.��(L�8�l�j�(�N�d��{�
(��w���o���F"�^j�z�Z�p&��}��"�A�:D�f����'��@�Ov�J`N� M�4�q#��I��Sv��H��9�haA�;7a2҂��`�׿})����1�h&t�إm#a��áI�Z��+�\�iu�j�cv,e���#Ge��my)oC�4M%~�U,Y���ĭ`�Y���X���8��5��;�;ݲ�c-��2�?�Ǥ���oL�p�mc3�R�£��k�IK�k�2c.�=#�u��w��f�']:Y(�f{Z[�4*MY�:KI4~�ť��dJ�]�ܹԉ�B���T�l>��taP `���ku���j���̒C`*sա]�{W��r{0�o>atȌ��8����,�ӰM�qE-x5�4�,���Ն5�^y"���.�����2�i�h��Gb�g�C��þ��E�6$��6��`�'�ƥ�	)����I�]�_�h4m�ƫS����A�7��}���6�\n�@cqۿ,���YQ��m\����"�a��X�Ε��N��F� l���/M�~���/k���命$`�Q�@lRi��kp�Y�4 M'R�@��Y�D!�ZB�d	�Nc�b�;a��������[��� ��7��vf�>8R�sD�)�|��]f��T%��DW�e-H����� V3T[`���ܟ�t�-�@ds�O�9o8�SY�'�|M��	g���X���h���Xb�s{sgg�kC8�-r�Z�a��~TU�7��*0=[{w<�x}��廌h4ApP�p�W�I��n~;i?ks��P;�&A�f$rz�Au�Et�y�%�����K�N�}}��v��Q���}��p�O򱄍�\c��A'��v�H(�kA�}�j(d��[�~����9U`o���%;� �׿8�L���3ߔ�J|;����Dm�@�ƞ��P�n��I�=S�8���[2,�s���-;A �d�H��5�=(��2�Ԅ�������m�A��Q��4���q��l��bb��EP�b��PY��?®}��=���UW�H�Z�	,&��[ 5A0Wt�������	Kw�PR�OJK���`'��Ɛ�ԡ�¹м�:�g��K���ws��.O��#�A��~ې)��p�̯�降V!!�d�5�����AT�ڮ@ ������e���q�a��l޾"�oJg�8E:��'o�M`E��X�t+��&K]�(.;�T%"{�=Q�h�\�����d]�`T󆗕�|M�z��e�aB����j�#quN���nK��$��V�q���BBd���S7ϴˁ{����,��=��Lɯ�7]�W�����R�#m'jcK��ө�ς=7[t��#Lbe��9/Őz�*v�C3Lf��z�N<�Xe������@�\�$��Oh$@���1�'cCJL�q8��f��~}hJ:�7Mܞ�;�lb��~�4fЊJ,���My��4Kv���iÉO��qH�����K�F�Ik'\��ç�+��*�x=౭���m�".�#����!&�&�9 ��ֵ�9GQ�?��e)m>��X�˽Z;������VnУFc��  [ ��U�$�ʈ$c���g��m�P�)��
�@�� "Nz�_����� ��Zh��w�/m�x�a|Fy�D:y݆��bM��\uHQ�>��-��A>��٥`P�zL!c��T&��K�v7�x`Ь�QͮC���=BZ�&����*��&�,U�,�[X�Jr.�܅�8�	j�	��ӳ�� [�U'��Qx
�'�u;�v���*��v�6������#ȌRXf�&sFW2�����c���+I�记���������R�O�:�N6�:�l�*d"�l���:C6���N���K/�����"k����˱�**��Uѓf%�Y�Th���:�B=[����K�����;����Xl�B��e����<�^O��a��x��z��� WL���̎"�JM��g3�֐���^�4���Yy��Þr�8��Ⳬ�<$��+{B`G7<����*�L�0-