�v�h��'˱����B��0s����r1��f/W���q^�q�r�����/�)�C&�gL��5�]j�G,�wu�I?�}A������'Y�n���a��"����)�� ��������CEu	E�,����z@��V�L�=c&�R��u�=��Z�^��)�L�d��ΚW��ܛ
I�q賚,9w(T����:��T*6`�z7x����H�
��v�I��O�3��3 �[��@>H���[Na��dC��*7q�/�������\���BS�6�2�[��"��H���c�e_sy&S�� �,4s�P����|m�썿��Y��MQ��Vn�ܛjb����o�x�]��S"H���Z��~H%ƈ�9�f�f�5;��t1^��E������!��B����IP��g$�j�%��!
���>�@�L4���-�E��1�����))>z\9V�6�ڎR�W�R�R��<�B��˪ɽ�S
�fi�۷�z/�;�����2���������?��|.f����i>XC��!�`v&���F���ܼ���Q�x���۫�&��=sF/2v"��B!����/n���d��<���5w�7�]@��,�6��쵳���;:����1ª����M���R�݀�q�j�ﳌ$/�I��j���HOj^�x�)�!�d���3�RZ�Y!]z+�h�jd�5|	q���(˗9m������d|����_)	���u�xWIh�4D���������c�>����(�����6��&�>S�T�a�jp�'�����$�`�F� }  ��D�xc���aBi�2�](���Kk�V��B]��B��AC�$3��u'�<=>��J� QWb�G�(A`�j�g��^JI�`��:���-�`�Vݏ�
�{�(�IC��R�؊�':b� MP��^ٸ:pF���_Ҙ�#��ǵ��
xs�F���*=8
��S:�t�9v�y\�������8��t$��d�xw����e�[�X\�g���@7�ȍ�@��b�"����������32��y6�J�	<)O�����):H����7��+���2��7[�k0�!FE!�4!u���d	 ���)�ۥ2 �~y�"�$�>:*u��V6����"ǉ���.�M6�o��H}�F�xہ�	���p�s����4`DeB�X�72�����['�L~���K_5�}�'P~�s3��R#�X�%��+�ux�P7���,�\[�<�(��\���id�<�N���u1�(��Z�G<���]��6�����;١1�E�ik*��1�H��.o������:�T2��b��?�bs[�Vz�u!Ğ)sH5�VbD7\����$���ע2L(�,;�c��8�ʨ?��P|U<
&���umI��{}Ͼ�U�ȃ�Cqc�`����إv��^+ҷB�Pq��v�D0V#�F��^i�.��V�ؾ��9!�P�Nn�!�ICƀ�X���Y�ޝd��bH�w^~F^8�dHٻ,��O���h������:#
�}�ĠO���#�nV�,�ԛ���@�pM��;u5x�5$�W)k����I5��9�9�, �(쭃�b&�`]��4�g��%6�l�@ck�����WF�g��1��Vv���K:[P!"G�f�m>0=x;��A*�7���X�4�L�����a�7�5���C8����
�/���Z�ḀЕ����trY�bi84l�4s�RIO_���!����q-kD���Mo���B�#҈���>�9G�
�)ޮY�7T�ܺE��������Τ�h?^t��Y�^��֚Ć�|VV�J^�Z�+����i�>��&�n������Ey��[� %bz�8�dm*	�C1T���D��,�jM4ɪu�{��X+�~%�}�a�NR1~�C� B� ��\��'�03t/6���a�Ĝ6�t_��m��&Js+J�y�ܡ)E�\h
�{�{�f�y���^T�C�#'7��k����B��ŭ #��3&�
�����7�dX�#�3����J����V����1ޘ��{�rخ���:�vo+����R���-�+6����o�A<�?�w/�Z/�R/��z��#{͊�w1��`�[��Q��E[%GX�}�������l�����N� r��e�|o����cKܷ�M���l����P�J译dlB�Mq]^.�o�����;C���P2>� ��$�5{���ͮyR�T����E@�~�h_�=�Y�<2��A�@�Kl��k��o�
X΀����u�W�W�~�&x������ܻ���(<�*)�d��L#s�"��IC��S<