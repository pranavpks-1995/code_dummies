|#.�b[��$p�N{ ��Y2SY��φ~d�%���S����&Ŗ0�
�_��K~1Ƣ�2ך�܁�{�� �q֞����<���_?5<j��d=!m�x_ ��.*Qw�<�;@My|��VC�7��;L��_�A_�_
cX{�.���{
��v��[)t=R�3�ߒ��ۅ>�I	K�� �|]���=��?���KE��m�`��ӗ  �B�����C|Q������O�����j�T�]�N��=�z�q�zf���đ��G���i������H{O�Pey�c����$�Dk�.���S,@�"�q�w��X�t�ޯ���50�n���pdRQ�������o�EK\���KG���& eՃ�$E�Nn���.?�ȉ�2TlI��� �J�Eo��|�Z�+o���{�Q������S栗�A+cW��b��G��1�VgV%�֯Y@s�t��o��t�	����
lu�"�P۾Z��$@ì�v��G�����XSaҕ���6������(i�0��	ֳ���=�x��'QU\M��w�76�岑E�Kk��a1�����_6Х�G(�_V�&�e@��>� �(9��^$�����j�\|�*����mQ���TA�I&b�i�y�t��W���b}�	�Q��ܝ�?6�����s3�rx0�`*A��֏� ���V,bz���^:#���ef���$�R\Tb��_h �|�z_c0�r6d����;�r������eL�p���h>��DiJ�U33����h�!�	��$�.�T�?n�[�&����.\6��*q������i���GM��g�A�8q_�4�2��s� N˹�6�>��"0�W����㯫�f:����:����̒peQA,�`�v(���a�l}�6�h��-�B��Zo[�`�7���X�y�Gݟ-�o��"{���-�:;[0��Lc�@�qD��E�@�{��߅ϑ,�8k��>�:QY�1��)_��j=��^��b�酯�}R)�'����]:D>��v���s��Uc܍p��P�-�(�Iw0��01�@�� ]Ńk	-k�� 8�&��9`�c	�l�ԥF鉣�ܸ�g���,�D�.���ͺ��:��kdXU-�{j�c���&�ހ��J�n�`�@�޹IYP3��c�Z�گa��u�ɉ�V��ŠJ���K3]]OJ���Z%i
[��J�����`�T��	� �t�u��<�㛝�@��I@�x�\놪!�Gcj��/|G<&�E*������r:�6�3�"u�����v�i�� G�ɣ�]���b�xᬰl�꺏���X�uG�g2ACqdjι��y��ۚ��"�zKa^9���a��;
��+�9>��A}X��fF:�F��8c�V��L������F�9��QЋ�p��"�!��	Xƃ[Gx/-V؏��|��������������n�P��5*�X�y��*�;w�Y���h~����l�p����������XY�
i<��N�F�,�,o�n�����(�3���ͅK�Vk@zo���{ǫ�H�>�"���>��2#��I�|�頲}6C��Jޔ��	E�J3��+#ɑ�/���BSr+Fnj7�i޷"�R?=�>\Ȕ��j0�R�`N�Uu�cԮ#�V�������%���7���^)�78�h�G���^2��p;#����DH�&�R{~)�w��Yz�s�j1T�Ww~� o��"Sip�]������@��T6zW�H;z��{B;"tWIp�����	߼4�� �vQ�G�'2E�H?�ܨU;���J߱l?T�$�Γ����2��:1Rgڔ�4��k�m
,f���K�lk^�QKI��)}2a�=��Y�E~P;��L�!�Asan�.���i���Ra �G�UP������Ԇ<��C][�V��>�Ke#~��dU:أ�;���s�#jl}3�I�I^�2���W