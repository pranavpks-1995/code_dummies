1�]z,M0�" g:�H,����6�H�UC)U��)4�� ƀ�h�`!��^~����H�!`R� 9{b�@?t�e/��(�) ����q�:WJg��PlKM ^��qSY9� �t@�llW �l�v U�90ᱭ����fL�c�[�)�5R/h�[���M�9ے齯q$1�G�xT�<J����Y2�UT)U�m�3���T�U��mϠ !�Z\Z}� �c���wx��`��`yV�5,c*9�շ%] YK���ds�K�4���0��O<찌��o���:܌�PT�Q���( �
O�
��J��	�y0�>t���o��Vاy�
 \���$���V����-�����	�&X�uU��R�+�!.��I��!���Iٍ�p �Xl�<   d�P�U��C��E��1|��{�,*Fy��j�?q�����O=�i�9�.N�9^4�� ���9��Ǳφ�3����Ydu�;EByU�a���XJ��<Jv	`kw�������Y(���\�P�VH�����Ӏu�[q/w����>�$�3��Pc�g��z.�a�f���z
+�%�I�
���Zv�k�$ �u�u@ҩo�jV�-ж6t�6��4�qƽA�hB���1��]E����u��7������zp�EPd������N�+хl}&����I;�9� ���,�fDm@����N�ïv�"M���+O��/�S
��EM���x,�fx���-MͲ�ł�bR�E��H��A��}��� i#�ZN�`3�-^!ob-��-��ds��-���-7ӂ��B�W�4ɝ}��꽆D���_.x6DT�LVr&Xhc��