33�DZ�W�:�l���4^z��>�ևJ�c��F�>�n@�*)�S=�&�q�N��.V�#(�S�a���,K���+���h��/Z�Ϩ&])������4�ܥ�c�%ҷ��2��*k�dr�׀�D���   � �-����A#�эN8V���Ӏ��K��-K@�� 'Z'�Ô�ҫ�b�vd,�#4+��������U��&m�ݩ5H� Hc�H�Mhtg��8�^��h�M�m�|�higs���p`'�S_��,�k�TN������F���Ba���x�y�]�M�|~L�t/�����|E��rM��%��J���xբ�(�K���A�����B����МG�� �+nTz�L#*���v/&mp vd�5���K�~栒��q�ɑ�,>aM#��6;����cfw����ZNwM��K�!@�58o��.*� �VIe������
�G(9j\�v4ByԪ��2B[ɿ?�;[�.l �����c>��_d�>D��'���H��������Y���G�v�flϠ�~Q��	���+N#ɾ�!E;��ߑ�6z��c��+ٝ��Y+�i�5����|�ZUOO0����X������1!5TN��
�!���Ѥ�%�R��F���	�~�����N�@�H_3M�U�7$'�{3�]-1S��e����W��\� k��c2Yv��4�c=T����<�(�DіG1���o%6�ㅍ���cDx�[�c� D߭ p�?��bY�Y�j