!WT�qP`����  <m<���U��������9A�-p�)
o�oɒ���g%@���4T
���
M���?��9������I�u��p*R�@0%�u��)e{s
b����XC�؅+��E�� �1r  x�{x.��#�)u�9ҍ���     !��������#5�f,�V���%��Z"�S��mbxMw�Z���x��:���G�z�e�'9
�gbp��H�wS
 m�n:='�X��E�6(����S��A�W|�Ir$ *������)ሂ�&ȡ�;�[JD��<�HBwR��V}�0 !���£0�"4�����f����z/����G}�j���:��v�o��I��$O,�������j�֙�6�k'F��	�<<��(*,e�8u�_ E�%���C���]ݽ�PO��<����i�����%x�5�&�!���[� B�
�v��  �!��Ą��n�#�"  ]� "~ʤq���=�U5�Y��ţ�������B�2����Lۄ��ra��^kq�p&�n���{��SS�L(NF1y�."�k�D@$ߎ6�oښ�H\���a@�Pߔ����M�g�3vW��D�fy8�L�o������A�T@3�0�k�ļ0 >5   �!�"�C���(	�i4T(3��ˡ� 9;�!F�Z���d�6��|������v(�$�������T�3��,�{f���pȧ��W|����L��0��IN,�n����h��������Ǿ�\ЗA8 &��L@U�F��C�HW]ܱ�y>  !�
"�d���B+���1 @  d`MA��ڵE�k�>\T�-d�Rł$A��>5K�D�w�����K�hRnN�ϮW$#����͙�+������B�u��?�J` V��@a�� ���=?m�� a���:m�r�pX	P�  ��+pf���٤/	����  ��P��   wӐ�UW�C����i6ԈsQn�� �s4��˒��R��1|^�k�N�:��k�@��Ρ.Zv�EZzf�,!�ﱷ��?G!��S�K,	��&Q�*��?`����ē�������%����12�s���U�'�����c\��gY$�7�$���3^�~�?/^���8�?��퇊�!Y0��
��!o���nĶ�l����h#/�2mL�/1֢̇Q��uL1y�<|YFd�W�TE�U��ʐ��f�c�����iDui��D*	2f�H�Qok�ơp����K�w�1��ɣ����$p�o�>k�o*��u�zm��f�i!��P���3?�
�d�Ý)��}�<?��T��:��B��t�35��Y��}~�6i��vF���T��XT�.fn���5����c�C�v�1r�9i9�״dn�����,�e��z6��IŤ~5�ZN��� Y8]^Y�Բ�}��uo'R͆�Yង��{�]�%��P0���H���;V&�œ�BD4@p�C�`G��##N(�ڗ�ޑ�a홐k���[zNy%4�=H����K(u�3���L����S�O��b�M��+�� �1��b�|Q���A�]��CQ��z�f��
�7�r�0�C=s��@P
6��g�Uu�5jMg4씥2�K�pOԝ�μ��q�}�vC���&.k.%�٩�_���.�Z@o�G��`��ڏ
��/S��X§�M;���XBEZ��k3Paqm�r�n�7"	M�b���(�l+�����;E^��-�j���� ��i�2xQ!��l�~�S��W����#������e(��?�J"S�Y#I6a��)�|�ެT�Pinqh�d��F�_/�%z���B�R�ࣝ�WU5V�}������%R�!~�֢G������ T���u*~s��<�')�)�i�糠�J��,��6��8Ա�wt|��s����9"����e����b8M�u�,�"�����|k���d*�(��x�{�����F�\ť!��{��.]hr� l7#v��c�ɘ���}p����m�/L�,�#��1��,3�5�U6*ӫO��(�����˙:�w�}��jB91���@?�l;悈� /K4�Y���)J����2JyTd��R쓈E�u5��3X!�{|#��I���������Ė�5iͤe��R'd��h�]��!JJ���/"F� ��\���3��bJ�;��3y�E4�O���UC21b�ţ�^�YpR����zb�=�Ҹ����H����ٳH�󨤰����-��� #G0�D��3ǴLr�+!#󠤇qsύ�d԰m�g@�۾\�|���*�p����?`V7��E�^ ��(����>-�h���0o<
�&Z�[���TJy���*9���1�0�0W^��!�'�1�e�aͥ�Êu�Բ���c��M��S	A������:�c�r$s��9%���w�@��,A3+!���Iݹ����0�[d�����w瘹�N~�d�Oo	&� �z|�l����Y�Z����DP|VVG^�����"�f�3엁�Q �=R��Y�4w����wv����׃�NWX��������wP�1E��3�Go�3��lO����{qʪ��qA�>�V�y�YL���T7:��{���Sǭa�('�JߎT��㌄Il�{A�+����E�.�u�+�E�����-��6��)̀�nӉ�18��b�mM�<��,d�|9�ϕ͚�1M�V��'�}l���V�րMY��X�g�x]l�U�HE&虌�}]�S���l=�n�$c4D*�b�AG�<�"�"P�]�+����ar6s}�w'��-�q+���/��m������{�d^v�����A
���!~	�u��&-P�ձRy�އ��Qd1�_T����^�YQR>��\�_��v*��8�Ƈ��&0����ys�EEx��s�UR#	�|+�}��)��7�z�'T�B�u{�JC�w��ƾ��Yk�˱�F�4���5,��Q���2���>���(��}	S,ӫ3�0h�TC6��W������;�Y���p���?��9J����ي�����$�V����YIoh'���
���ꮍIJ��㢽�~��V\Y�ʅ�0�˿Nx9	��,��b�-2�D���_ڜ�m��|��q?v�,���R���:�Z���i�A�@�4��>�Q�m�ʩG�p��N;��Dς ��0�u��,U�e"����@Qq]L<�ĴH=4����f[biq��G�N`-%�ޡd!t��y�����v�+��˧���i�^�K�V�>���.H�����*�n#�>�e Ӑ[��T{�+4T�����,�:�9�u�iK�0���o�rWo�,֭k�5}��Шf5t�qW�7�(,�NP�4`p���y1�j����~�^�V�8
�@�@������4������^�v���P9��<�_ ����e/Na�����oS�5��/<A����i��e[A|a�dȋa�HA1���#W�x���i�e��w�}ž7��o��%[��?��/�_�F&j~I�}A�=��Z�f`���YI�beo��x�M#���-�]HS�7�Z��"�C&��ɯ{��p�Et���o4֓n�S5�e�`�4�l@�9���V�M)b8�f"h����,��i,{�.�]0\t��DF>t]�&�Vw=睓������ú���ʣ�
\��MIJVf�P��ץ�'9I҇	>�[s�̓i>�L�tT��d��������p�Ë"�[�/��yO��U}�}��}(|9��1i[��̆b[�czj��FnW���uO�5�J�tF��y�hD	���7P��7|�ǱEӰ��F����v����n"�9Ǜ�"���tz�56HI��x��eK�����xF��h���k	2����> 0s�A��|��υkG��͙�K0D| �zq�|5�G�W�f����F���Y+N}}7��o�uF��+>s�zWؐ(S@���'Jxu�N��jXzr�.����h���݁,B1�s��x���]�xh9�U���XG��f�oc2J/�Q���M|������-'沙�3!�s@�L0�� |į�)��-��j�5	y�9����E4����,gz�,��|T���.u�`2G��=�We&"��x�� k����`�!���}�vT�.c?�Y�.����k����h�����{��&j/�a��/����h�^�T�S�]��\�x:��!�b�L8�WT�+>�]{7b��ЇM�`��3d�� L�C�n�����j��-I�:=��3_���y5�����zx:+sk_�.��+X�i����DOe�!hS��!�GTF�"�&3������wo�6}�Wj�
D�É����}��|~!��G���0!DM{�n���E�f"�U����部:�����4��T����P�(L���hG7���ѻy7�kߕ%��l�k��'2-�רM�<���ۼ
=L��S����Jf���@J��h�Q�������̛�M
4ď�#�r?�u~��
�_z���W�O�� Q4!l���RX����� #�SaٜE�4�������RoJP�ҧ9�WLͥ���i�����X�5���t)�8�8�O�6�i(ԛwy�b&e|_���NL)�m����VԶ�H� `<ոw���E;T����$�&�ȣN�̠��I8���o�Եơ�����@�W8׌J��h���0���iüA�T���Eg�>��	� %�f��QkoD�Cc��i�t0��fr
�{ƪ��U�z�� ��:��C��!�F�TX�ˢ*�n�ARɁ�eKw?mK��>��	-�e�I��+��1�=ނn�Ƶ��L
ƨ�T%}��G�$�]lxsy�
_�
"�/��O� �k�n�����П#%�`��w�2*6�{yC�A��R���$��E'E�K���W���r�(�5`�� ��HA���P1�����'{+�ӳۦ�m"|(#e�����*ՋP>�c[L�	:�Ӟ1�;u�P��A@=XLfk�+�����i�g�_��S�
m�ck�Y��~�����k��Ȟ>��^>>���ȱ��� +��X�Px{��@;jk葬*��	O��.����>Q!���_6 ���!��x{hH�J��  

�%RW�c���$�YV����Hs�K��J]�A����_Ȁz�#�u��ݳ�y*�'���&�&B+����
B�@D�&yF�T��:SrQ��|�e��;@n��FNY#B9�9����-<M������%\��6&�:?8��E�ݮ��?֡o���9������Z��=2��H���=��C�N�1�4�D ����N��,���T+d�[�$�V�k>��y����@;�]B�r�]���(/���J��H�W�\�{mo��[��fZЍ׌��v�?A�1e��?exad�1�N�x|���bi4<�;[_'VY³fl���T��M�Y�Y��mB���0��*7]`rƘ�M�<�����#Ǒ��Zp���4=I��\��C��[aՀ�ԡ�rT��9�J��}��K���Z�<��I0���Ҭ�j��������M�d(�D�I�k}3�!����W.:lu���s^�����\f8N���W!�����yt�d_� �eAh��r�<L�
���-j���뼕���ĝZ��./#�g���� �o�����֊��B��!T|� ��q'T1f��ju[������&��Y�D0��[?WLu:0�&U��w���b�=�0
��mp�0i��@9q�}|�52,��NIe|��������L@+�X���nTPg����m%L�����X�Ɂ�q]�)�f��~�����	0Y=Z�Ǜ(�Qh���Y���!"���%�j�W��q��~����rI*ø|�S@;��	%#+I���Z�"�)�����P-)��iF�8u'���K_�ޗ+���b�xwW@�$DCj"4����d��q�m�JE4���C�?���ƨ)�J��d ��d�XW�7�EP�:�Z�\��(�>37�h��M�����2��Mc���W0z�x��)5�^6��G�GG@~6�/��A
�)�QӾ�#Ie��Un��UYӨ[�r-�4�H��=�~��~%�חqlC1o_+�4��Z�^mD�LL&#��fz�lz����pQ���zZ��	��l�61�H}��Aͅ��a�Ӓ�	�)[�s,#cÎ�#C���|w>k�mt�����5��}΋��콬�s�ީF�8S�O�Բ/�9ke댃a� V�%�[����4
j�����Ώ��L�Öu{��7���|fG����9���r�����-��Z2��p�����V��	�85��,f�'�!%�O�ݞ�R�}�v��� �)&��rh������_(:���
�Va��<?I3].ʄ���4ٍ��5�.&�<ʁ��`t���&�u5sA���J�w���@�NgO@��z�����\�{c������쇇yj���3�9�|��gF?^?��>Qh7��կ���W�ܸ�(\[a������D��_7�a?{������9������'}���<	��XݑC��ɠL��<�`�: ��lB,�+����hJ37�{!g�+���fv�j6Ɵ#/���v+�i�3�0Ξ�A�~t������*]���?�8�W߻C�2��s��=AQ�"����?���Zi�� ��O5.����L�m�]�ђ���7a�W(�k]�*i�4�-+�`7TV�ƹR��R��<n�6V��0�� 0���gB�Av�w�+�-�#$ͥe�;	�zЀ<K�	3dB��%݊Y��Pua�.�o�Mʣ@Ճ\8�w����lJ I[b{���~�y�C�,
6��jj �ȝ7����������$�m&^��Q'r��&A��GE/.f`�M�n!���zY���y��j����{�f�bY���W�Q���&���S�w�>�1���~�� o���4���n����9��̾�p P�����W0x�I_�ND����{-�o�QO�,v����9����T�Zoy�B��#�����N�&}:��C
�5�����>�p�ꛣ�;�Jr�HH�-ѓ�&R�Z�Po�G�"�� ���0&��"�-Ӷ;��q�������o�TH�`��[7R,*U�(����9�!��	�4w	���l�ۙ�TxN�!k8Wh��f�v�� �3���ab�w�@R%��>S�p!.{W��cH∢X״�Q�����R�|�KS�)�ф�ު�j����|WG���N{�`@f����ޅwl��~��@o/���9��3�������7m.�Qb8�PP�JϽ�V��5�Xw�ݭ�����q]�f��CM�֖:|*(Sh|�����C)�Ŷ��b�������t`S#��vU�U�v�$�h��_g|��q��8�^ޥS�_���<���f�� �o�5�� � 5ֹ^Y���e��=1�B��AH���c�+�3�!nAE�襋��.Ls����̒��.��6��N>�;p�v2<q�tٍȲl�G�F�Қ�I�궿�Ƹg$���L2$�^[|��tkz���Ԗ�ȂuWQ�}h����Ħ��v��3�XrI�3I{���-s���W�I�&͉Gԝ�-yHأF�u   �����,t`�1P1(��oh��E�	���"��W���k�!;!���Z����M��	T
��c���D5Lif���o�(T�d��ȳ�N� ��Q�'�~x$��<w������ШǦ���y�^�z�~�6���ZR�"��۟�H]��ٟ��]�d�ZS�e����*�9q�bT����sk�?bR���ν���p�>7���w�����oX�S��ք�P8�g�{������"5|��a�L��Xk�VY�H;�h4��:<&�ϸ��� ~	��ge�b*-����as�$�8&����?�T�G�@[n�:��'��h�q� .� �<��f�.�U`��\ 꿅N+�Z�A�Gv�ˬ;uD��![Aϒ��׊��wYM|�r��zex����j[�'��\D!�2)�9����ԝc�XC�]������vBzwO������@@�� Ā�^>��~֢K�DӴ�Lf�Aucv&��">�i�oWi�20��6R1n�<��A��#��=��eQl�ռ�*<�s��� =��Э�o�"�R���'ۣ��m®�Y�kVDYnVp��Ł7�bW�G����{''F�5l;B�(��.{�`3�[9-�� �J-Q�`��I���}�X{�9�ʝ�?m�ĸ�B���%B�5hO9/��i���`k}2O��{b���A�"��/�t�QN֩������qB<�D
���G'���Ѵ���s\'#s�n~�0j���
e?�ֳ����B�uyr�cw�D����'fc�8�� � ����鹱V�0d�E�
<�����25��8z]kNM�)�e�"'����ݩ���W�!=H��2�en�$��DG�F"KN��E���F=oa��tl��`�1�;`�f �� V�E!8�澆�&��ێ)��d�r'�7T(G��5���w׊Q� ��׹S��,�'d,�%K��L��hU2����V^�Vz�Hy����/�r��'Ċ��U�]�{bHg����/+H�U�uG�e�!����֏n�N�\�L�/�c����O��v��Py�M�]QM�b���p�fW|bkv
q� �_�%ԋ�_ٗ�L*[<\������
&Se���*���'����q��Wn�m`9ڠ\��q�� H?��u��s,�>��}@�����u�Wm�2O.h�����O�����5��oFpe���km�y�W��