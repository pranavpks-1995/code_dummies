t2��2��U�^�U�V���f��)�� (�W딓�jM��
/�"�#�_���:.ճI9<�Waq@�߫���r�[��B�
ܱ�I%�(�4���Ư"�f�z�|��Az�%E3��wI���4#��Ym#����:�����u�P�ȹ&�]�1ɗ�5�>݌!��JL�B���z��{���԰�T�)��.W����U�tnKs�1�`��'pbW�Y���6�3��}�>�-�0$�8�w����/έTO�.�����^*�&�{jh�����
���	r�m��6���	WPp8��O9�b�)�?�>�MP�$gKB���q��Rs��le[]�O����h�j��:�ndb��	�=��/d	u����`���h GE��<�؜ޱr��N���Α�T����l!u�57�1���\ɯF� �����ṹ a��'��;0�̱��h�������l%��L(��=9M%��Ͷ��	��Dj�,Mg�}�e�$k��HPd�#��4Kכ=�d37��y��R�Z^U��QʫhF��ZGeq�o��B��q\d�����!5I�a>/7��A�i��V���߽��<8<"_h��,�g8F���t\9�{?�c.���ڑkB�-�L�,����r���V��^��RP1��3뻘��_�央�Xz����$�D<A�ܧ��ʝ�
�� ��6:ѰR��B����uL�;�q�|Wr����A�G��ةBo�B���X��o�ܴ�����#�/��v�N���B�庎�DS���55%ʍ|�Ц=���տ
�6o@���"5�����Xm��\J\� �Zd	S�˿��[�q��!_�m��f#B�w�k��S�l>���2t��C�q�׻����s���J,;����>��Z����(276q��_�mJ�"�f#��o g��}ۚ�D�7���j8:p�WI�͎��Cԓ����~s[>�ۃp\$��[�K�5�|4�K|��O�h�Hb[�6M��\C"�{>�aUGj��X:�pk|2�LQ�Ƕ$'J��2��W����i�s�㟯я,��K�y�0��[Sk��%o���c��
lf/b�%�-��uW!�י���&���C0���p�v�A��c.�����ik/5��hr����~���{fX�rB��e4�8�Щ�~���	cFDY��a7`�r����i0�:�́@���	�$���>�K <�\�X2 ���ն�1L�r��Y�����n�u�Pr֗se`��9TA�SH^���x����wa�dĄЮ=��������o�O�uΣ�/�2�H\���\cY�X�"{�0Z�b��f"�h�2�pjK�EjS�/�f<����!����Q�n��x`voJ���Ƣgz�Y͞����4��`�\%�Z$P�w��l�_a���e}�т��ѹ�a�]DI	7�F����q�npv�!�����Ȧ�2�B�³����d��H�j�������Ж������k���*0\�}$rmk�o[$�<!�1q�&�Tr��Y��h3Qa( ��ϴ� xp�e<�}�8�B� l����a��&��.�Kc1>�j�`�F�Le��v�<�w�@�Z�+� ڝ�$7�~D?����J�����3AK�&CG�w��AK��|��f�6Όǟ����<��&'�6� ��7��� ��KG��Zcr����P�m�^��b�pn�/Q�����>ֱ�� ���x�<tҋE�曣o�����K '%�qA3J`c���p`�<'y��R:�y�:Т�l���9�Q����yd:d���Y�ϖ!��Obk����]̌/ǖ�{��Ok��!�`�� ���ad`?���ORJ�H�=O���t�_"�[-J$	�����p���,#W���i�5Vd�iQ�ى
� �~A�S�J�I�-?�?�t���(�Ь���覐��?��Io#�'���b��F���,�M��^��P6J�2� �1��ۻ+V���A��m8�tF>J\�w��F#�	�ݓ�T�	0Q�ft�l�<$@?�f}��^?�eQ'���4n��	f��(T��$�������>�zd@�O�Aƿ�0�.˥��\��G�f�+��%\�}�E�r��?��f��aY�k��v�yA��иC�Џ&@���e�z��Wx�7��4w�x،6������q���2k��:�y/��l�7�Y�3�/,��jF����~~ы�#���,�u"�*�u0�:O�5o�p���%ɟ��6��/-6@c�C���Y�f��փ��3��i4d�rF�����h�^'Z�N��ac�2���K�]��
53Ա�W��"�h����<���!@�w�V	evF���T����}�V{ ne�`��g�<���:�gyiX��bD�2�w$B���sR��&gOoV�_w����<�Us��ڑ��h���WJ92��� ��Oa��y�	}2s򘼡)�G���61�[�3�*�?������䪦P������͖s��qzr���$��-���v-���ag�c�Bݥrˎ���S�v
+t�5*q `��̓�H�eÛ�A�NƆ����&U �֛!BR�$]��(ҎAh�Ϝ�X&
v��m����7�
����3���� 9�"/\�����>3{�W4z�����{���ڮ�ַ��� y�`.����	�S]zX�JǈXS��S]t.gD����d��%��kn�I�!���6κ��0��W�2��	���xn1i�ב2j�G�m�%
w�� V�f�_�D����[��  �!A��4�\�C���  ��"%R��c�tY���!��R������R�QE^X1ǝ�ʺ�^|����c\��������o�ε�A[�Tv,Y} ��צA�-�+(G6u���4�8d͓[�>�66�,,��LZj��ZW8�Qd��(̕�*CF��.��rpɸ�=�و�����,a�@f$��h�˿u]����Fy,X$�s04�s#�|�k9��Z��<k
��Tʪ��s��T���E/��䙊mդ\��`��=Ϣ����o���Ϭ���rd����	�`�Âw�����3�1qP�F�<Y�S�+@]���
0Le�(Op���K>�t�0Pg( �?~"��Ȥ���p]uA�$qy�t�c��y���M%�3k�8��ө6��� �w���@�L4u�����������p��v�D,߄�7����N@��F0][�Ad����}�}(�TO�͏�9NWJ^����Ph&��-o�ݓ�r�H���1��n�.��>`"᥂�Q���VI1J��Zrk`O9ܴ�;�����s�Y-����Big��3V�ŵ��>�%�33����&4>O���:Ow4���NA�鞱#&����!]*��HV9��[klN�B!��lO��,��i�2,?��-R�Ͻd�0���޿�sQ3b =k���9ͺ��G��^�m��:/���N���17/����҃ɚb���M�Hx��h)l����j��� �O��l������4�k]L�i:`�%:yzQ�+��g]5|~���B]