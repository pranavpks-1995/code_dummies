�{:�x���G�KzhT*|�������A*��0w{�c<�:)��s�����ME���Ř��*�>ɢ`�{��
�@�M�����T�*�*��.9�� VRf�8rTzr���I��E�+�47%Z3��6`T{U����ۙ�8���`���9�d�P��x��GB�!��4W�H�%�0x������z�A��P�y�Z|�4� r	��	�:'����v�߄"�[6�#�����[�3��WgW���yb��--q�rEnn[L�9����<��>�2ھV9���p�;�"o���Qz��o�jk�����B�����d��+��}@1%�|��?��;9(3�0xA���=�� ��At�ʌ@��6¥���mVo�{�5���`��	��)nX_�C�I��c����^����Tht���~�5��l���j�IGЛX?I�b��_��;�g�Ц�W��a"�N'�}�׀K�d���ERu�8г��Rj����V���f����l/��êoWe9&xr�j�$�����)�q�E��`�{}>"�h�A�A�FЫ���n���Q;�J�;^'5v�f!-J��=�}o�?��ҟ�*�����B^i�UB���h����Ԇt��x�dS!����
a��x_�W��L�8 � �{@���NpvWEZR��r*�=�(���l\"������E��A� �$�H�8k=�Y
5��|ac����~ϋ��B�ˊ���1y5�(^�Ҁe�B���bb�|���j."@v����6��H�i"q4\{J4�֢�_ՠp�zzN<V���Z��!�Ӆ#�'���0�P�ˋxD���u�w�b\h��t(�v�Z��}k��o�r�z@��J�>4���	1}�Q�]�݀�
�V_��>p�yh���/7hg�����
�?�`~Kr�3�!���;��<��BwP�f�7�T�/��⚷^�y˶Zm��	n�E�`�By���D!Q����d�UNZ�.�[��L��AB������fu&�!E��=IJ{��\�%ai�^��ȒPK���Ԗ�}��	1���?�S3���7��������;<c�"�a�)h���b���V��1S�1��I����\x[ӿR�@�w����mjrp��!��\��=�if�i3w�g�ʬ�T�%A���)Y�����j�=�=[Mv��E��w��/�L�����p�f��o�b��4���c��Q�/{��ݛ�ȡ����I��&�����Wg�li��y*˴ZN���n�ʈ`�Ί��h���ӆ_K���S���o�m:��72
6���(���+0��4�r��1�f?�u�c0ە���'�\�r�!�,�"�9�~����{SC�t��%XhAa�d#�RC<SRx&׏��F���­I�ѣ�&�C:G�j	T�4�n�����v��'6j�s�2��:��T�eU�u)�b�������c�q",֯��k�Ak���I�y�>>�f㤕W?��|�'p��ca`^t�l�t;'��+�|q?�}�2z9~M5??�NZ��
�tМ���d���h]������n�{�1�Ú��IUR t�k��^m;�**�˅�3��9oT<J~��ȝ�I{������2љ�/�4�X7a6R5[�r?	x��[���l.����`�VI�O�����`M�������>�6�ī�B�:�,����V��{�rA����T�r�
�f	�!��Ɇ�1R�uC�>�T6҈��X�Б=O���@��7�]j�et�֣�����Ю�x���6�?�:�K1u�Ad����Oڎڨ �Kh?��ݤ���ٿ���E���	�<'[Aք'=n�Vܧz/���A��/�#���X>S���Jq}zn���-H�[�f�(VU�Φ�yt2H� W���R�g&���m�GH�e�H�wU��"٧@֍K[;��Zz����,C�'�d�}()Ӣ����}kkYO�wBz;�U�믎��lD�lp���,q�� ��}쩄b�ٵY���g=E@���4�l�Y�0��Y�i�5`�1^q4?�̮UV�2�={�p*�'�@�O@�E�*)х���VN�*�f�;�At���W� ,�;ć:^�b	H|5}���7���)�}i{h�HR	��*Ť
�?U
�p�"j�P3R#\XΚI�?�L=�� }4�p�����rXЅ�y��p�٣����K��a��I�U��v=E�߼B\�K>�7+J9�%�w��X��EM�s 	蚛w�[_z9�ؑ�G�i��}+�\���Q��C��Ø(�Y%(%^��c���{�%8i�r���=5P��W��g�ƒ�h�Uy�3N��O��l��ԁ*���q1i�S
�;U������<���E�!�\�-�(39�9Kl|�6,�%����[,&���Vyn#�I��r���ԃH����~ôY]�G4�-��]��Ψ�f^��ܓ��s�xj8�%$�6�����ۑ���mXz"�L��� �<I+�p��!%�A��r����P��*�Ŀrn�R0�C��>P��¦�2�*���qg㔏f<�j�9b�IQo��������T�7��B���z���`8��g��%�����n2��U���f��Pͫ��-��?`��au�$�j�u}�B��x?�y�?.�9X*���EL��6�~p548���}Dp��_�k�8���%�*U?��"y�~��;m��p��Ё_*#xIr�=}��k���^�d����/�����3x��~�\����39���-�?��^�o�3+�Ҿ J�o��p`���v;0�m����&�
A�Ѽ=��-O��S_��S�N�|��p���D��U�P��PC�(�G�m���Ƌ'��K�g��I5lbu�.���Nz,q�e�_p�9.%'��g؋�������umyP�IZ:�,�,IA@�6������]O�N �6��e���)��m������=W����CZ8�B�D2W�1�ת��[0r�AL+ӏ�a�2?�6��g��O���}{�O��n��|^�tzv>XQ����?kO��PA� ��k�4d+\�>L�[���ZI�A�w˲A�hi��?�nX�m��7\c�)������A����.�e9f�h#�2�@���φ�͊O���d+��_S[��A>�#h�0 Q/���&bݍ,?���W���\��ϭ��8��U�-|~l��N���bw�/	 ����T��@�f(���o?��e���ʿjS��llmD��QA����:��2�>q��S�69��އKl{�$oi���~HҨ��pjB�S���z�k����o������@�O��H�^a�c�:�������`
�d�)�EZˢCh2Z�^_�lf