z@�L���]#{������(�\��sc�����¾ {�N��v���	�%���c�&iِ)�>U=�����M~��DH[L�=JRr�nޢn�C6&���ܝY�I>4�}W�����.]��K�.(NM� e�:�T����N�8�x�ɀ߸N��u3������;_���[�
�J	�p�X3�@r>��O �ʍ���[�5_��4{�G]�?q.o�6�r]%�D'7�z&�'z�K�j(�P�"S�.f�J��1��bO��V��ǧ&C�_�v��R��ټ<(�?�Î�"��l�u�kSNMr ����I����Bm�zA%xO$��Y4�)�X�B��3J�J�+
����$Ð�i�(�x?�2��=�1�J\l��;�μ�Z�����w>N�ss�3�>s
�7�h�����֒д�ʍ��Y*3Mt���������,�o�c����R��%��2Y��]ƽc���ې�5��<�U���;�tE���k҈�l�4��D3ǝ�<�v�x�uE@?�
�B{m�B@�1"<f�wqچI|UW�{��z�j����K��<��a�7�5o��n���X�p�}
�>lW�q�L{Ԃgh��eLr��o~�M�f�$'��{"��1� �	���o6h{A����TNi����f,WY���)�}l����S��t1� C�ƌ>,ƫ�� TУ�~�	١�ӏ����;�^��uO�M�ed�ڬrU!;<�ͻfl,r�=��5Cѫv��_��1�< �#!M�^c��ӷ`f�-���oq�����f�"?3�b��c�F�L�e)I���`��4��i ���#Z	[� <��'U]��'U�3ͩ�<y��=~${�B[N����#6
#��f���ȼu+l)����'��U�Z��ru�틎���]�D�Ö�q��U~����V_����8''Ƒ�����.(@�C���Ƽ�iN��f����#�\��77�OK)#bl�@��o�0�3���T�q��^cQM�'x����Vsr�j�6X\k��� YS��(�v�P�걂;�.I��f�g�������N�;l�a�i���p�����,�ƈq�Wa��E҈�
e�{�P5�>	<�\�ڪ��ލ��MZe�2'��sm��!x%$�񦨘Fq�IΫ�!Xl-�tc�u%��l�2aDW^}�^e�6��:��>�C�sX�p/��e��xJ��\����� )�	AxS�P�� �������Ѡ~U�K�8xP�hJ�΋�J/ѰX
��l�������F����|B�8�
��>ok^^`��A�\�����d�H�7�ќ7+�����
;VC�m;�������U��@�PK�H����H�S��	]�cb"1��U�if
˘9`���P�jk��}����=�%�ٓ��yI�9ML�)/B��W���}kW$��!�Mt?����=�M����?����e��%*��aM��ǰ��qr\��4V�;o��~����[���1p�������q/#�c��X��]:�������&����v�G_�.�Vq��bZ���o�-0�Յ���c�KslE`�|���?�kg�c
��z���=@qY�����۵�J�2��R��
���$�v��j�	�WK��gj�?�^�����wit�?j��w����bN�_��m��vx0��}h�*zw��;��́V�V�vV�k�M�Y�]�@�b�wWi�,��*�h���7�V��[�Q���#N�p*h�J3��sL��MuFJ�.�F͒q(,�$�л&'�__j�Nj`:��*�x��Ơ���?��%Ht�ZCwrx�b`C�C�O��
AH�ѓVڗLH3����:2�j	�A-������ݥ���N�G��Q�
-�u��s䘡�c	p(�ِA�`&��0u��V��C�l�S�1|JJ0���ѸD���&N!���5���X6uKd��G�D���,�zgVL����I.�v���>��2*\�ɷ�/G+:ג��%���1�2Do��'�Ps�_��J{Ne>prhR�(jl:?/9��*�K�ɶ�d���}�� jt�?�G�pj�'"���
�p_�[�<�&��.w�`�h_.�l�~2�*�����"��Z>�;8��wJ8�r/�^E�C�(�R|�Xn�}
K H��W�b4�t�� ���ϒ��\ ��N�Ug]v��:)��������%�:8����ֻ;C��D@��D�Obշݔ$Oo���n{���ӕ�=i'm�����[�w��e<��2C��9�����۰Ќc�%F/L�ġe��v��k��`Qr�Ƥf�JY��\� ą��%Hѧ�9HH7�y8���\�xTeѽ:�GS�3���_���=+��#�����j9���Oe�`�9���9 �X	
Q�,�MTQf?g�+��?ѓZAƙ���zizɂ�`�W���A������ѫ���t��$n�2/�����Ʊ��zj�f������`ꂷ)���v|�z���it�^���)�)[��x�خA�����,%7-yH�)]��2ڱe!���b~`٫ �TsK����o�\C��^]P$�@Bz�-��h%�(�G�;�)c�R�vAq�G���B �0�ۂ��_� �ȴܞ����Y�~�50iS�x�ٿB�:��BU%+���*���y�b\���T�n�49iEY�f���C�qot#ܚɩ���ߡe-L4j0����]�`zI��f���$���kB�B�w�Af"��$7���s���4�:�t��'��Mj���S�b�cSOQ�Ӱ-��sR8q��h���U��ƌ#md:w�{��7ǎ�U1{in_�<ƖF���q���!d5�]��
�i�6.]�[Ƒ'�xP�h�^�^�bA�*���Ї�r���2�s����vt���M����嵫>pq�p�%���,�r�;���
F���N�oY�m�"߅[������h]��ը'rƏ��� $�mE
�1r! ���WǕ����(*���ܰ����G��E��	  ���%R��c��ؤ�zqDT3���g��BN�Y��\��UC�����*�Xgw%s�r���x`QR�_S 5I�p����`��G����co�] r����)�[��nP50�?��E�|��Y�c<3�{N�'{��Ǥ�{�o]�� ���j�[jgI���E+�U���W��CS�q�w��x��W{�-�Dl�Յhq[����/���>����*���\�ω=����P���~��&�U�8��;]}e�������\r�R��h�W��e �j�c7�b����^;<>s�|F���
�����o��S�ͥ{���Z9���k==�]�3�*��y��ř.�� .��P"��;�O��p�^N-D�_�:��}�A�U�2�<��R|�����Smc�Tȼ�;�pa{Olϓ�t��\iU��۝�?+��qޅ�i!�V�PM�<YK��:n�����X�l	�����Ӹ�����"������Z��(_���	^Ʉ�z(g�T;V��I�|+�i!+�|mA�.������d*,�'͎���Y*ef��̝@�r��n�'Լ[������w�wU 
\��]L:�p��!
��D���i��sy��ʹ��L%NOF���3rW>�(���>Id��]L�tٙ@WKNٓ
�O;/��1��c����U��P�R�N)En?Y�&��HK) �1z���g������[M|w$�"y��@�n�ľ��v�l_���(�|?�CyE|��A#}���r)S!����Y��Lȯdľ��4>v�j)�)}�e�+���|gWc��[4�m�u� f�u{2��8P�"&*�g!�o�}J$�\&�7J{�������~���tS�
YSbi�d̿�0������5���%*W������,�+��?���|��0��b3`�pU��F�v�w�3�N������ߓ�
-�ո�QOCz�5��(ܲ�w��Y���n-�D!M_ӭ��ѯ�g�P��S�S�'�9G�7��Oz�J�@�|Q�: �q�����y/�����7��O�G�1�%s`����c�NX�k�V�֋iE�-�mf)<C/N��7-�"c�ұv��(�'��Q�$\�#���0�ժ�-�5(b;"Ca�l�&��-*w5�ɁH;���d���[ˈ ��{��MBmwoW�9�&�%�A<��%���A�H*���x���!��W�r#3�Ĝ��?���Q��4��%�o��s��p�9`n�hl
��Kݎ�'~y׍�Q\���y��^��*�H���ɝJV��R�jؚ�B�v�վmvS���3 5��͕�	;4�@݅���uQ9��/鎛lh��Lp�@ON5�h����
���~���RyȀ��pJj��:�5���PhM]���L�}���!��9�
��y��U�4O�TitI�i*f�t�B5��  - �����,t`�ԡ"s#�q�e���A��E�9l���CcA엫HV_��>H���[����k���,�V��U���C���+|�(�r)�g}��� �C����<݄+�r:�4�/c�V�0w|}9�S��q�'�K��#�N3����( ��n1��Ĵ�:�U���C ���"`.}��w�Og����%nj��W�3;�:2��J��� �G��d�D��Z�`@�50@F ��U�R�Z��L�_�*�P�� �(_�}��|�@Ho��2T���E�s��L��!\D)P�`�K�V�/)[嚦�;���g�_�Y;�%����'�l]%��Q�-���n��t}�eJ����\�B���|��#�>�C���l��h���=�����D3���s>�2�^{ 1��d��.�,��6OO	��Ĉݿ����>�+��>� ��cm�y���-W�9�|���uq�+��5��q4&}�-OJ�Ё�|�"����;��A5��|y�� b�;�����v�gXK�xO�LW~�U9?/��+0'`�Bf�2   ^ ��-W���H�%GF��ã�p��[gQ1��Hw�4l���&m��^�g4�(T�g�S��MRhe�[�t�{��b#�}�z#+bG��M?�f�t�H��ph�5z���¨O����$���s�@��'�/�lu7R�O��ݲ��G��E�Ű�p_�Z��!�p«�ٱ��|vi|�����BA�xm5q��Q���jn.���BΦ��U&�(8-)�N�c�,��T�J���.�i2_[(W�=��@Q�tE�"�h^�Ft6�'4�84����i]L9.du�)��8 7�7L��1F�����q f���-�9	F+���ݞA�Tp�џm�}gm�a�-\i�φ#N����yt[���b�K1�W��e�&3��|��=s�<'�I��v\z`�@���� �E�ފ�����%_���H�J2�h�O�X�}@��~٩c�1��|��@�kE����2]q�ɤ�
��i���%n�߀��MU�Z>�r� F�p�II���t}.���o��T�_,8�;�M�����~�w�o�9đ��s*���h���8'�l�4!��a��R�Ώn�f:���Բ���X�E]��©�����!�����2��:�` E��vm�>x��@R�>�v��<]!�bV�N�y!=�w�Ӳ]�SI=���)�O�K�
�#E�b&T�){Nf4'�!H�6����u:,F�@� ����
-ĀD�%��I(�&$ʐa�UK��	��<���d���P�	�"p�%�q K�.P���@��aUI�׹ʉ4ݺ"Le�-� @�!��?���6a� Y[� �},���2�3E�o�q;4��Y�ǐ���2�����"6��AZ�A�{�w�`	�](B'|�1 pS��"�  4
N@3նG�K��>���O��gj@�� <��ō"���� F2#�qj���n���� ��Ph!��VF7��FB�U >�.2�6��*�M+N�`u}oo� �cu��u����;�]X���w64�~=M�O%��e�o� �Zӝ�N5� I���@( ր=�x�/�T���ZD9:m%p��+@'\@Zn*�� 	y.ܰ٤*�Bc�)D �!��=)@�&@��f,�������6�j�S4��F��R�H�V�G<�����*�&�r�ӥ�![]U�7��\���7B��l����������r�� �" Y��I�E�,���0� ht/���x�Ҽ�^EX6߆��`V�c��R�d�� -0�U$$�* 0  8!��-� #v� ,��BWa��4�6��t���e�
oa
F���?eos��I�y*DRdŖT��4�D��8�M*S'���&��Z�0d����IAQ q@D�@� 9�����'�U_Å	q��r|{x+"�?�&
s� `�!uH���   !��P�(!�A���ീ����(�ˁ��a��텾�-C�[ԑ$��#rDa�7�+���bz5�����	^u�
M�G�0�++�����X��O��"C��h�)$ŠP p, +��؏����\$hWH�V��t����O��mc^����5*�  !��L�!k��4V� �Sp��@J�:� W2��:�R ��E�A��~��C)˕I78{�g;Q�Xa�4whF�=|����C;�(1���0>�C�βIB��Z�*�D�`AB �@[�Շ��J���t���)���
^����R�
�  !��A*A�@ ��X �>��>cR��R*�)�Zi���Ʃ�!��/bҡ��C��r�)�DUV�����(�A�3[5Md���{�Ʈ�mܴs�>���?RSŐ��|��&�@����5� @ 5_{ɔ�2�����.� ~� ,��S���4�)�(��U$ ��(0  8�S��-   ��h��W�C��j�LC�CQn��~����t�׮`����U��Y{f�"ǋ��:U���Yb��0Ն�5���Ĕ�p)�.��8����P�C�H6�f@l���#���Չ��㚰�;����m,{iF1�\�r�4�U���������7��D�B��뙱@l���SrפB��緐�Ok�⭆�EB��r&DN\�z��z��[�/���:��w�;{��%�Mϱ%�
u�r��zB��p�&Օ�yjZ΁����<���
WƖ���*MIs�j�Q�iu'P���w��#�zҊO'ne����C&O�E���JG]u��{�#�Bc A���zP�f����i�Lب' O"�e��3<���!�i�Lܯ��YV�8~t��d,�ֺ�{w��ӿ��3���X�'B�a�z�M�����O��E�t7y�j��d ���A\�k��d�<������i!n���3���9��#�o��3�N�xI\Fbd6#�@Ү{�G�}���c�ݎ�pj�|�g�\��[�l�p)�[��4�P�%� =9X���q_���z�=�S/��([�@͙#���4;ج~Hta5p���<��*��i�0��R X}�@ͱ�^
�e�nr��}]ie��@���B
q�U�^zފ�s�_�lM���1����UF�턚�����IizE/��~�@ENvܵS�C�^І�@��ݦ'F���mb��D��ɷ�$_N��q��E"�.@�R��-{I�Z,=K�v� �5�h�`�>늊�k3��pt�� �
	Q��a-޺�oFx/ �>�K�-��HN)y��C0{I��o���t �haJj�"�C���]�Կ� �v��k>h՞���L��@q<��sp?��=ݜ�Pr�'�.YIu�7H6�j���3;1�svxW��5�O__Q�*��w�"��-����tʗr��9T3ɔ_(��'����`�w��O�����a��Λ����� 
Y��"a�l`% pN�'Lǒ����:g&��`}z��lB���;I�Eq��s��2JnF��^�]���F�ة"x�(��+�f��2�c�{c�(�c(���vQ�4�`p׃�f�,F(�x���tPs�$k&q��`�K��c�\,���E����'5�ϲ�ݙ�Zx�y���b�A�dn[E�E���9���,��r:@I�jt�]���{�A+%ſ��y<�@hT.ÒN��n&!�-��[�2m��%e����@�3?��S���ļ�f/X�>�ps�I�m���0�5�-�9�w���Zx���Ĕg�'y@�Ŭ�-��>h��jK�.��Ty?��A�9�_f]�a|?BC��a���a�BG`�_���E�4:#��>��x�Ď������@��g��V�4���M6<�������I󠡣�+z���gy�6G��� �	b�}�u�q�`��5c+�JRHVk���j>���I��ݧ�g�?7�,�(�>�:uK9ڂ��޸}�ѿ@]L̾��R��%ׄe�k�u�X��k�a��;	g�.�+=k���%cEB�&���B� Q�m�}�x�@�ok�A���/ X�7<�j_8�E�7��n)T�[�c���5��M�z)�y��샑����b�f7���?��