/xK)D�) .����em�S5���� ��r�����M`���;ӻ�ů@r��3�V�F��a)J�����mA���"$hi��:�A�|G��s�R��{Dp桡."�{�����3@��c����������w�54����*��dϿpi�ц��x�;f���z=��k��$�������7�e�	a�a������Nh<:����pD�������ʓ��:]+�����tI�*�ŉ��� ��KZ���B`��`��І��A�m�M) |�>j&��4�g��r�ȉIa�|̆b"�o������s��̠[��-�?
W��h�6?�Fo�)����Q��?��"�T�d��@��D����ZP�c��\��	2}��uw�¿�8�5r�Q�
�HM��9��̆��t�c8�<�j�۴&�X���0UDo�n�NEVL���,b�9�C�88�e,U/,d,�/�i`������l���ɘ�S�
J$ԅh��']67��9| ��cVb2,��'"�nV}#�zCy��ua����\B��leǘ�g^G�3&8=%����	�KP������9�E�f�PT��Z��Ky_�����Ԧ���ۡ�N��^�q/W�N�m	�ɮ7��y)�y���Ϲz�V��{������f�/������xug���[�	���E��d�|m�>�����!�И���@`h�D��Hd�)�ʥ+^�@b/"@��M�h���i�+o�we~+�]�L@3i����AA]I��Y�L��� ��U�(r��+_#�+9Ss^GT�����������ԋ��"�ЀZ���=�~��e�������^
�K6]�ۇ�;��/L�+6�T��	�b�ⓚD1&��:6��J�}q^UB�/�[BG�J�b?h ��� ����T�V�����!�$��FH:P������x2�.ttT��!u����X�3m�y���R�W�<�d"�p�56)�^%-��n4��kavv���c;�,Kx�����4KQG8w˚i%�J�NJ�x���H'~ղiW���$/����^X�oۨ���-��󟵄0:꺽�`�T��
,eNb����
�@y@�������?s��£T2(h+�\�w�\s�B$؇1)� ��1�?��<��.�p���/��:9�X"�T��h���X�8���t�T�s".ȸ&*�E������(�FXX t��*[j�h�Ĥ��<b~�2���<"���P3��ºvv��l�ez�p����4���LK��� �č��}�9�o�աK��)��`�bvW)m'Y��Ro��p�ƻ��6@�_y��G��D+)�j�]�ǔ[�7
�á�؅�@�����a��0��k\��;��P�~9�ׁU1�����F2x4&+0�线��%ӯ�q�D�F�t��Qh�hI9ʨX-��{�v��rO�\o���σ1����L1�}�������f." ����p幊�OH�b*������vG4�L;�4�PٙSyx�<� �2�:i�fE>�^��k�r���Jҷ���m% �V޴�'t�Y�4�Kgz*�u�"E�!$Ơ��M�o�Nq��es-�\ÃzS����ii�1�QMjq����O�t�K��]�����o�ǔ�C��_�P�FV6µT�N������s�z{6�^�Y�v�><q���$����G�k�݌=h��z���#W��������Xa�C�[���'���:��?��[&�������NU�3�Q�5>!m�2���6W��sQLT
9`0'+�9��|w��-w���lCb���U9�i6���#�-�����#"u3t�[~��~��Ǜ� �æ������"��5Oί1�tf�Eb=��~�č\�UuH�����]�������L��9 �?�5Z���8n�\o���DB�� TT�aEi�D_z�`bZ}�wA!�R�4C�E Sh;_������3�aP�z�0~{��NFk�����v��'4MT��7F.P�|��%Oػ�(�u�:��㫾�x�O�C����kB�쿹���;R�beT1��ub&L�ўa$M�gbG��*��2�-V鐘 M��S�)�b$K-��Թ�DگC^����3�R��Kr�U�Vo����<���_�=su�@@*ݷ�t�UHe�؄�6m @E�<FJ��c��d�B�_U�7 +��bw?=� ��-���Ѭ�*A^��hܐ�{|�[�Dk���pΰ���6�����T�7�ӽ	��A*�ԇ��&�6�`�M���B��_�C����p�(~�^�T�j�r�%0�S��M0ƶ�fr���
����Z��U)Q�z�RS�p�ɝ�͟�ݙ���4�<b��|A��1��	����ƴ�V��M�@>Ax5SΛ5�l�
i
k�d�S(@� =i�{γ��8(#V�6�w�?V����.)ؒx���5G0���+��3~�Z�� n`\��gP�[>7A� �h7J4^�\邊��aH�,���Z���G� ]��z���;p`���䆦�8�.�#�S����g�m�=��b�\W�#���^�8,C;U%��+[<b�W����s�1�2jQ��~D_cy��C�:����~Rp�8�g��}J#�LB��*۶"��v��z�l?�AW�x)�,��3���֩�w
1�L͒��U�����f�ԲI*X��P%�-�F51��;ߟ�Äa>���{3,��I�,F"w�B�J���K�b2@�Q-%i�Yo��,�����׹�YQn����U��	�h��E�`WG�@����A�A�y�~
�#�y��˪=y�djKg��WE�U�g ���������j)Tў\�iO��n��[[��b��8^b$�I��7���\3K�j��;��K-�A����A-	�?��LE�	���vh%;�� Q���vL�4��@Z���_E�ۜ�K��+�u��
P����<���Gq����mN��l�����*�t'��A�j����QuHf��ө�Gx�
�  p�'R��c���S���նZYe��<jN�:&ؠ*�#�|�%���I	�r
T3�^0��`������`(�&ΘJ�%U��<2\�rQk�@�z�)�_�K���LK�A�SyR����r�|�F�)���U���j�{t<�T���������N��[b���	�3{9qPX��͖u�Xw��b����=rn+0������Yk|v�p[���������t��b�.�b�/��f#+8���T׷](��P\{t��e���P��s|���	�����29m):E��~%���ީ�R���6�+ ����������e�c�j U㙟!�I���s�*q�ۉ��˾KY��콫��w��}���j��aq�����XwX�D