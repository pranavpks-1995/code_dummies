u<"���f�I��1T��^�Ɣ6�ޢ��vUQd�����>����"M�伸��Ԝ��{�������kh�����[��>Ѣ6q{SZ�/KC�#	����M�m�L;��%BF�i�+^"��mHfb��$?�]��Sdv}������W����Ǘ�4D(dS
%���P�PE�	~:ȸ1%S��!���B$��+�iXEIUoH;�v���,d�fԎ�q	cw�j�k�OK�VWk�Aw�eIw@�#�kL���J�L��_-�B�0mDɨ���P�s c�I�s�����y�I�,g)-�-�7�9�^,:~�M�|-M�k�w�o@��dF��N�s�ܲeuO�0���B��P��8Y�8�s��������芟N�*Eq	#�Л�������ϛy��6<���:P���3�<a3;@8�H�*�z����#��������)���
�{���{S�����,�tٜ�ʲ�d��j~����ن�-�ߴ&v��)+"3���?��:��3l�J	Ͱ\��c��"�9�"�5�1����S���+���'@%R� ���Z�D��%^vIZ���d.5������uZ�樧�#@�3��wJD8�U��SdD��a���P�*qPA@��J�:���M���t�((����U�횥)���x��� [>X���z�mc?���K�s�V|�\�_����]�zk�)0嬱�<����q�j�안W7N;��I��|�(�4vͪX�N�3��_�+l.O�c��g����]k���̖�T֛� XQ�Y�R�ws�V���x}�`������?P�z�O[Va��@�h�D�B�[�ť���ł#D���Nվ[D��S��M��
����؊�?�L������SSP��Zo�ޮIFlO�z�p�H��Ɲ���r*�9��h;*Æ��`?��t����}���,�-z+X�و�̈́������y��k*��� ��g�H�Ӊ��̰��
�N�Y�)��2���[�� �A�@�o\T��~�@(���g�i*<&c���D��4(hi�؏��7z�T7�����_�����s����e8FY�f�@V�du8]g� :�[6`�"����{뱞�2c�C��,��k�1`�%�H]uy}_��OL&
9%�
�K�����}%������h"�P��~��U1{D3NKC�GN�wV.n��V��Y^�]$M��H�kڔ������(��n�(�=J���Q�
����"���zDгUN��zT