nW�A)��  ! ����,ta�Dx�8��eX征��g����l���W+j�M���kS��^��^<�� ��y	5ii�\�r��-Ym�3��rLN��Q�7�Pmv���D�d����/���`O��z�ر��Ћ���oh��UJּA�]�i=�;	��]/ͫ`�X,8��P=qy� �*�O��M���L��b�g��r�j�71K��Uk�3r�=G�QqcA ��W�+�2J��-x�q�������[���wE�y����% ^�pT��Dp�����g��NܣA4�+   , ��-W���F{��I%�jp�we:w^�>�e�.�ֺ.n���LL������Zf�^ċJS甒�˝03a�i�`D�M��n��%1�f��]U��@�c��:*��	ϕ)�Y]�`}߳#�����ˑ�� �H�X�nV96�,������h�s-=����$�h���s��KF����q[�/:��@����S�l��H��0���y>��F�� �O/V$��1�G����:W{��C���Oaz�;��	��v�3�e����T&�L�M�o����q���VI��X�p�c���