^���V�Ͳ��}�B��1� CX�W�CTkK�<
�GW�rF	�LRΒ�Ve�&��������C؉���jc��ℚ���sm���-�AY��O����x9����&>|C�IٴR�/��8A�?�R���WJ���;�O2���zv���W��f8��w�N�`%ބ���q���ב(���()b�A�!��b�x��ɢ���d��
XFɪ|}��'���o��z�7e֞G�δU���$�VtH�n�
�)4tVf��g���h��-�Y�eG�&dKA��{w4�i�i�p��?ʑ�~��96�ׁ�&T�\������"w�����!�1�i��11*7qk	�jS�*^Ӧ,���t���:��y7-d%>UθT�����Euv+�*���^`+Ӆ�RX40n��-ݚ���`6�\��I"�����Q��Rb�$`)�����-&���9o���,��]:E��N%ǖ�Y�R�%_Pg(3c�|�!�36k�}!s^8?
:l��)�	�?��6��~ �s�X��l ٕ/Jǯ
�s���cn�D�4Y��qx���w"��RaF��ŉ���R�Z�@�c�S0{�+�����˗��g��n[�\u�1�-��]a*R�=�"�T���A������	S�o��OVfFO";3����`O�ZrNJJ�(��k�^�	u/ܰ7ƶs��9q�?�q��Ă�yr�Z��罨��M�Yv�yv�Fu_bn"�
�� 6��C!0��bZ�a;��L���;�r(a�	f�.4)>�sn��&U�G�Sڗk�����7 �S�w
Ua�֕�;��ZtK��?��MG^�żGِ�Ap��;X肽M���ۆ?��|�Rb ��(�����Ԧl���F$�}�k^��M@!6�Ƕ��4N#J�X+�[4�ϳ��{ǂ��[���h�@&�Lj.	k�s��+u]�4e���;�w����a�($��n,*9s�(�qM��G�3Y�;,�[J[ �'@�{���n�A���zk��j^�Aꟁ�������#6�b��A@�ˬ���:ԆؓÓhߑ���[��r��:��Bb�  Z ��U�#��0�TdX "�Y�-���GbX;�ԉ&�K�7�b���ȡwW�|���g;�;N\�w^���-���y쬪�]
�"2W���Q�w�G`g���;S5��� �	J0A���{zƙpB��_��|�|*k,_ym{X��RS4Y��"'��3G(Р������d��A��%��\���qx�}��ó �e{z2.��8�D
W�����dC���s��{�+�`�	�Hs'��m@���ǀ�?	OT�Rע��8��������n�OO�E��_K)n��]����ۗȐ�ɷ��A�9���չ����L�2Ј�e=�Z��x�"���@u��5`b-�iv���"/���v�u�.P��a}���]P>w���!xB#Vi{��R��i�~��$/�A�rBJbD�H��X���·���^$�Z�,�h�~Jt*b �8���3f�{�`�a����NkX�FVN8���30���՜7����ڇ^΁#An�����Kv[�=(����.İ��/��Z`qD�^q���K.�kh�j/�h��Q�D�i�&���/����QJ��5Z��,�<����'�	��X�Bā1   � ��u�&n���P�t@R#��Uy�Ŵ��D-Y��P