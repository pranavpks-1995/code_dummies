>٦
۳:��R�簹�ٯ���&�է{�AnN��]B˝��6�0��76�Δ#�t�MR�7N��g" Zظ��q#*فe��B��ֱ�T;nl�x
�������u������6����8f���{�rs����eJ8;�Oޕ1���k�^2�M*�XM%�5����CiƅO�n1�FB$QtS�ޒ�<)���I.P��s���ց�v�6������:J�q���}	�ù���X*�˗�A��1���-<+0���G~F�y"��BXR��*��:�r�[��w�{8z��XMNͼ6���B>�L�����$A����d�{��io�����ˊ���'Gl���5h �/Z����8>b[�1��`NRp4��K�N��b������%cR�|?��Sf�j��ٔ��'Em��S���$/1�J�؛Q��1��>Ț=��N�����V�2��	��-_���	޳q]H� ԯD�a'b�Is���~����Ht+;����O�T����pBC�B�2���'�5�?�nY���g�>���Qg���n"b��'폦z�+���4h�s|= �Cʁ	�  ��'U_q��vH���p� ����3[=�p��W�3Ǜ�z^��Ki���F�=2n�`�D�Qr*3��W�{;��ؐ��^��tcV� ��Zɓ%c�kEv F(	ce��6JŘ��<�wÌ���m748��K��R7�
�ɴ�#^�g���)��K�]����ÇO��9�Ａad �sRDk�է@�y��G�Jaղ�;�;7��p,�y/��s[D�:��Mi�9�иZ�	Ƭڪh5���56qRC�&��Gi�p�#�3�v��Y�\�_�y��������$N-`:,��H�5..��A�Q�T�r�,fǇ�#�r��$(s���ݖ_e@W�pT�r��4�O��(�����
J�5(p��ΆK�I�Tq[E���I��o�W`�њg��lD+�D��?K�B8�;RbQJ1��r�ᵗX#;G4jvۚF��i��q�zM���!Kju�р~�>�1�����"H�āH��'ﵑ��bV	��I�������ꙇi�f���Y��Bq
���j8W;s�d�D,���tz�XE5I�IRD���HZW�(�J��}/���SXQ�i���Gi	�fx`g%���i��Di�
ez[7��=���d��k�J�l'�k��ؽ�uG��ٖ.~�-�wo�Zth<�F�~[��^���s����O
j�'FGZ�E�\T1g��È�g�`TY�g�����;[�hU�:����4�!�-��A��	qn�Z3Ib�O�����a�,N-�Ъ����q�"^����r����lJ�Js�i���[h����>)2*�R�I��@g嫛Ƀ���Q�-4��������������z�ٌ��鴤�ut���͈*�`F�����B��,�kƄUP�o���wè(B�G*�ȋ`�l�o}<����g	j�#��?�W� z�t�JW��_5�(>+�$�`6���B�	J   ���U}"�F�d��-Dq��6�E>��j��� {��W��P�T�H�,Ǘ�Z ��:�J9�\�W�X.j0�'��7���[�xtvN�����\\Y�%OW#n�� ��s�� ��V�J*ж��vmek���H�B��ѳ~&�8��M ��:��u]��]b�U����l���8���]p�#4\1�J�~���f%�}�M����Z�W3q�r��i�	p��ϕf���>4ɶ%�o%�?���*Y��.ժQ�^��z�º:���@��u��`�HF`�����D��KH��55-�fTw��/�������}��5tw~%@V�L8���jF��4�+��0�;��(��i싻y ��v6W�O&��Ⱦ�\���bX�R�@�_jQ���z�x��5�U`��̬�B~�H+�����sM۹~��icbvs�Č5��H)�pd[ߑ�s^Ӵ���E
�~�Q�v�#q>���Vǖ}b��+��E����/�d8��R��(����*=G�~8*{�L����ţBg�	s   _ ��ԝ}"�F�R\�L���P�"ㅬj0�wBM�W���������sb
����yAQI3�ґ�C$E�}�����˷�9w��9�%n���Su�T�����{\�1��22�}?Du`�H�A!��L}��X; �����h��O��H���)_G��_ky�t���9�N(��[	��) (-l�!�Z��g�/,����-�(�1S�-M&v����:k�[�V��MJ�|I�@�M :B`9~����sdh��OQ��HD6��Wߺ�p�Y� �����;��t�KS���@��:�.�i&{��3|8�rp��^�ns�C�,fb@��p��ɾ ���� G~���u�R:N#�����"�.���J�̈�H�9kco3��o���ߚ���y���@��0��V�Ddu' ����X�n-�37d�n�9O]-3ֲ�i�oѡx�>���]H8Ky�&.����#��E�哝�w1&������?~�*;�[Y����3#���~����6B���I�.�zE������dc����j䝄EݤR73KU$�.��?Ocʢ�9�B�hW�>s�y�dQ��C�w4�����IzK:�УA؁	�   � �"-���:0�ɚ2�������/������uzn� h{k�:���R��kp���xV@U�غ�Jzg����~�[��@���~�VM�`h��&�E��f.f���(@b���wj�ᴳ4.����Ĺ�S�dg�L��=���ty��K�!Ń�"N3g�a��y����Kg���؟�E6�̦Y2��6��iO�
�����|�ʫ�����$Rݱ_��[�s�/� �@%zo�]�K�u����]�W_�^�~�e�m�]�X�N��RbQ�ԇ�3����Iw�WT(�0Hpˠ�4~Ԇ�2�XB��4��������ۂ~�b�;�>7��9���3 ٦��pW�z��󨅂��4����D\ަ����A��������J�W\���~ӑ���~�ꍷY�O��x�M9��a��ڃ�ݤ�v�p<Uvh�����t��/�� *�!��(�ஞ�
�p�T�
�   ��0�U������Lm�E�B`�5���K��/
���] �����_̎8V?|^��u|�g�	�>�sȾӟI�݂�?K�n �y������`����}΍R_WhY��V�=A��s����8c����ژ�b��#z��[�U/��O�;R���t�:t�ML���xK��y�r��e�l����_�͚�_||�b�ϰO��*���ƶqB���U��(��ᾯJ� ��
��h��7W>P��t��[�,Q��Gq���:,��pdb��N��&��=�R����N4��7�� iWR�k%ަ%^��n��yO�/`�8
�?�� �%;�Ue_�3�0���a]��#���urV���_�-�䨿z��M�t�[�gm��w��� N���̧��r�[Ǌ�w�e��Z����RYFlP'��KiLd��C���"_3���o�2�c�}D/2XNǢ�w\�I{?�.����i��(&��������W��ނ�z�e����ߓ�p>�� �V��u��
�rXH�P��3q������M)<�y�cv��G�9Q3|���e{u�'�E>\�L�\Ύs�MQǆQ�x��@E��@o�ÈiuW�{����u&	(�+�}X���~U�@w>��n�tt�F��b����f�ۇ��n�Y���a�P��{.a�pDB��l����0:S%j���]&��š�rx���4;ޟ��#��b�pD�F(g�w/X�1��&����x8\j6<BM����>4$���z�	7��繢L�ґ=9֔b[cU��TD[/N�p���#�#J�T4A���}˕��iÁ�qDQCg%�`S�_ZJ/��Du�e��`Q\y0���I���LW��K@ULp��z`t�����k�k���7+��nM��(�*�%J�x>��\��<1��1�C���j���Z=K�Z$w�Q�[�~��R8�1ck�ì��c����?z��)y5�CF��q��)��~�?��c8���<-����}
ڮpǨ
y����7���� ��yy]��A���UE��WO���0M��:�*�#-/�@kȒ�PO�mV��V?��aK���]Wi��/�,e�����U�"W `50^$z�1R�ӄ������j��`-4Ӹ�r�Ay�C��i-Œ�Mǎ���L���K����o^�6m��f�JP�9�"3��Gr(� �7`��w)3�ۍ��'�a�P���o�p��4	�0�F��W'�Xp|{Õ�S�L4Dk���Ul�Q�Nbo�R���S��ucpG�E����&��9�UN�	������8LJ�{����Ugq^�śecQ0
��d���}!���=������)��!K�&��pCI���,*��PEE�Er>�uVW!��ǄZ�{^wO�>�����B�yj�	GB�`�@�'����uT�\ O!��}B�E!ɩD�d%���{����F�3��0���J���k�2B�HX$4�����V�og؀�*/ ��C���]�c+:k={�R������=�;�3������k��6sf���3�0L\a!s��3yÈ淯�d��YY2Il/���4�Ԏj��	��^!��" ו��9~�3o!g�= e̀�h2��ꓫ>��s�h��!}�F������Ƃ"Js��KY��᳝? 4>CA
S'��Aa�~O+9�%���p���,���@��͟��}$��x[M��C��V��ߘ�f ��e�=	�}r�lE�Do��W��{n8�$���$3lW����(�_.ј~!�kO�K�2��{'(6m ��un1����$E����w�t:g��t~��tɒ��J���U� �[�m�3����+�m:y�[���
ˤi)~�&��y��$�=�}��
��`�����br,@�sy��,�|0=�/�~b�r�t�27vt�i}��D�jm�>ЯG���~�
~^�[i':�q����	k���)fH|�nȝ��FFj�ق���2�h��ILx���=�6w堙S�y�	�,�FRn�0�g����&b���{�-2�d��U����W�I�pe��'����fs+Ų�2�}�Ix�X�i�;½�<���n2����:Cw�5��xc2d�дdY�;VZܵ&Vb��"[3X%�W��1<��~�J���M��ֺܝ)�<v=���\G\��Z�E��Y�M��A����u8�Iy�O�����ۜ��'p$"���y��RQC<�p�5�A������\���C����x�dg]a�z<W�Y�L^���GY��;�'���� R�r���=1�d���L�?R�%g�fYm�-�f8�,���/�4O�[�!K��i�v��Ri�
�q,(�EV.�Y֩ aL�x5��c��������3���N�?��Q�q�V�fd6���߅��2�U�"L��Ia��P�dO��̖¸j,C����+v�.�V����%+��>�X��?9�Y��B�`0G�=ږuhP�$���֣(���u*&��,#-cm�Vlbk��+S��	p�k`2.��4�6b�˽���za�!L���(˦�A�^8�"m��/��n1;�X�¦ߎ��
T�:{��y�®�)=Fǫ�ѱ~bl��h ����֭TQ�.��%�:īsk��O��߉XJ\��gV�qY��/���0qޣ��j4z5>_.9��j�kj�Ls����@�(}�����Bu�:���b�Y������D_�j��J;�kUZ�,�/	J�DV�|�5
˩�.SZ͍�����
�L���{X�&�eQB=�v*o9�w!�/�G���i��Z�'�HK�t����ƈ"OU�Gz�a��9�^���9X�Bi-��<�x&�jFzbL����HW��3��ae��FXG�,5��+�+������ӧ7g	���ވK�vC��?��4	�2����A��g���(4p?��ކ�X��du��u�a����H�aھ��! ��+�cM*��&�h�}Boy�Da���SF�]u�+=J{�����%��UE��y5�al��e�)1%���E|���4�ɼ�S��HEh�?Σg��XМ��v1�s�W�$>��gCV|of"φ���g�E�pl�r��cF�W�E_Q���������0�\ܑlŬ*�M�׺!��v7���ޠ5�tP�� �S�@��f�5Q��<>@��N+�`����G"q�5�H�{@�bh�it�}�j�s��e�&��dzaR�S{�2��H��Ͼ����Qj�		h���I�Tm���l�<��>������Sם2hC�^��w~�4�m���?��6���N�T&&�zC�/�)b��?�ݞ!/��z��ۈ�j�=�K���F�סj_��<�>8K��R�$�߈G;h�����r-������[��Y���q\^��"R<=�qi��K�O}��B�Æn��˛׹��'�jv~����޴]QǵW�8�r/R/�f�Jv�]{�w����ږ5�9K�
8y�񷞎����]�_�ۤ�4�P,6�E~��=a�����qkZ�&!�b}�h�f�<��5���>�a����Hߴ+��^��qk:3�j�"μ�@��ߏ�
h��rb�TB.��p)�s�_����o��ٕyh���8$3�qzHd,]�������C6�bʘsǖ��ᧆ���K��LwE��d���韾�O(Dk�F:�?5�@a�y��;�Z����W�@u�UvaO��!��"W	'�)+�4�N�6�p:�z����I:1a~��k�O�S�x��J	�������&N�AB�ex�ʯ,C	*"�.�y���.c�Lݓ�n��NF/,�V!�?��vlD��#_�֧�KK\ K\�h�⏅e�=���r�h�@�``77�S�A][�:v3�R��@V���>]����{����lRi�U����4��C�f��14g�5.ˎ������'y����7�bku1��n�b�P9X��&k������L�>oR��i�����K]�y�+��Q��H�UJ�������-����*���y�ړ"'�X�\$�h]+^��!��@��}ֺF�9�A/!&5�s�ߑItL�ݗ�x�R �_nq;s+;����W����->M= �aY�y�)���D������Y`�s"7��=�f�ռY=��Pv�v'�YW�V�ɎAܚ,��
R*��@��'a#��!;h�&�������,�U�ߎ���N�m@����m7FrU�?���&��\���)��g��>٠HR�1Yq�hgװ �kw�a.#�v�������B5��ӂ��a�&HX}�6y������\��;*:�8ݦ(b��2	LU"�?������z��O&�΀6��H�!�]� ��������zF�I�M㌤��`|����j-�iH[��G�N�Q�#z�ffO��u��B�T��/� ��z�;L�rVX��W��_��|O�<#�m��֜�v ?�E����&��,���r�P_���/d�2����{�Y��j�wY�|s�N�����i6�滏�O��`!��AL��4ل;=���8�Ѹ�1��ɐ4���(b���PL��ް�-����z$%����蟼�j�8ÂI�d�V��XGއ�̱��R~f$�FF�:FR@׮��9Rʓ�>;����n�9�ǎ'�f�+���0�b�q�>8͔P���64|��詳V���%�e2�׼Z� ��Q�w���7����i�첒��e� 7�2��٨���8��*Rq��g����ϐӴ_|G���!#h�X�Ǎ@�ϱ}*���<Ѹ�'��}@h��j,WK�g���=$��Y4�'F�����G��%c�K�ȸ���Nhp�T��ְ����V4�^���h��=Md�ɏ��k�c
�`���>zM�(��.?7����z�E�嗺��#�:y��u�M����i��㑗u��i��N��x��!�v]P����UWiG7�UG�m>ؓ�~K(�~f3,�N���c���T{kO��.�<�Ң��
C#��x��P?,����F�����0�N��b�^\�w\r����_y��fM}�e�5q ]����l{����Q������µn�G�|�(�x[����0�'q7?�ѳH^o�rm2'�8�ς�R��ܙ�Ί�A����6��z��1����c@�rp�����O%B>!{�$�Оo�$eE���Xl̄mp���6�zr�p{�č�4-^y���+[��yg��[�T���c�W!��<�U)ժ�����Z<���EA�
D  9��%W_q��'0����=0�`�q�ɒCW�ue����9YW9S���P�����1���Տ�%c rH�'��6� r��ə�]��2�-�x5P�e����$�
&�׋�h�~z�O���"��wt�q ,��ݡ�H��ܯP4��K8"� R
��p�Դ��c�e3ѭQ�w*����#�<]�-��kj���K�4g)��yP�Mf�l�ju,��2�-:���M��F|��fM����Ia�'r!_���V9�����瑗��Z0�wc��)�3 ��KN��W�C����9�R�;��̶�Z����n�z��6B؎�}F��+
8]-v���ή������g�᪳�O�4�n8��C�69�aQ�4�XH��S�έ��@���L�cʁa'���0���7��@�x��_��l��3��P,5�r�P�ں�����PҌ�"�#Г \��@�q���yK���dU��U3�~8N��#d����'��phQ���"������c�D"C�AA���lu3�+�?�K.)�3�����G���ȐJث��F/�f�*]@0_q�4�n#[ږ��₳����W �0���Ü��8t�߆��t�$a�xT��k$�p]��G2܆6T�S?� "	�Y��xJ�H����G8k���\>��b�Q�1��t��;L�DS���ID�T�B��o���3��_WET�\��x2aըj�*ζ�k�,Ν�D
g	��w�RTn�mp�2���80���%U��<Z��Y�|�L��Z2�B��c�!b����V����O1�d+�6��4��������Y(�å�fK�;����K@)���jp��stt�����d��i/,(�"�#4��7D�FM�z��(��� ׾�6W�<�^s��)I���q�0�U8�d5��������-��`�M�(��;��Dފ��5䕒��+��[�]�c��u�,����C:���W��t�i����T-�O��F��ezb ���������}N�=.�'�,�V����{(<��Z�9Ck� �Q��FoV��Ӱh! ޘ�=�4z��-[��/C�m��ߒ��b�Ngw',���-}R+Q0c V��4�T9���چZz�F	5�܆�K����w�)OWG�jyNF�A3+p���`��@4��`��ͪ��@�*��]�k'͸����Ή�ca�π,,v��|駾���?dՑ�xv���-a)�(og'qt�8s���Z�DA+?Qb��PYb���٪�=�m5�#l�t3���Ne�Цاj��@�u� '`<Q�̡$̥�rV����7p�[t[�0�A��
  � �f���,taוB:3�̟/�����^ާO _�SH��]��+�
�C�W|���H�E*���q�-�f#  Cͫ��}��n�n��J�l���{]¿6���M?~�E��N$dyC�����#PZ<a�s�Q2Y����G���t��G�L�����.=�������:S�jb3�E9qLO�����F=<¾|�w��[R�
�)���C�V��������TyK�j(7fx� ��o��B7��0����Xp�R/���۬x��0L�h��|� ��d~�LQV+��_ܑ�w�ST"4F  �	�t�FBcf���	,��E��~]W��чĔ#��l�P�M��xb�����j'Xh./cC������2#\�~�R�������X�%Y@�$�)-�+4�Z���w��H>�e����ߍ�ik�/�
�J��B��
n   | �-W����l�e��Jr���Tq�+�g�J. ��k�.���!�N�8%�1���0�cQs:��Z, Mv+-���'�_ zC�׵��Y��)��w^Bg��fϹ����X�* ��G�Dj�Si}���$qt�.���E�44��� A�p(}Ch�M
�j�����g��Y�`�Ǒ���\�#����JImS��e��H��  ��W�x]�����U�8��J��~���ݒ$ĥC{��`|���:�_Q�%�cp�Y���o�j|~sH�����mx�h�������^A�3�Sm��k������zTL�Ǩ�����þGb�bg�:Ó{e��/���r��R��A���x �_��/&�mQroZD⭀v��jQ�q/%U�ba�w���I��&��B�l�޶�x/���K�,PJ>G�]#��^���V�D\��U��p@_�� ����/]�����8j�z�iT�F�C2�2:,q*�K�  �.��'�4~�Fl۶ S5��Y:%�y�9��%&|D&���_
��\3:ƛu���k	 ��.w.Y���B����"��^H�*r_���+3��b�U%�
X�H	:���C��C-ʢ��w	�Ӻ����ټ���F�M�.y@�E�
���������!y�В�)bpc�ś�WE����x��g�w�|�y�����e��*$���P�� ��Z�7���eƊ��h�Es��D�����iT�����PϦh
9��f�Y��4�>�ֳ@ M�����Ht  N��)�%�U3o�|�^ߢm�S���H�     `!����b��( Wn���5�Jj�:� C-�}���W���0+ܿ;��Cep�]�s 9��C�Z�
,з�Ę wz�r�a']����{9u@D!�[x�S��A�~�?i|\�:~ҋ/�@ ea��	�Ppp(�x.�cw���RW��m�    !��	!@�b(��ڥX��:�1�HΞ��EʋӥG��<��g��/��(:.[���"��v�A9��gt�O[ߖd�`�۪\w�T���6G^�m>.���BbNw0^F�*/8�	�|���!)X~6�gy|@` �!���c��1 9x1*�w��Z֒���ț�L��x���z������^���b\�5Uĩ��z���e%��[ړ���D�j˧wxge�X���A���&�qMY��g����|��W�qG�7=y�Ο�d�Wj��@%С� o�0PN�!yLg�����(  !���C��*vL��wWk�:3A*Q&�{2�Q�q�۲���|>�6l�\n��X~5�Qg�"��������M�*+�����O����i�z� ��Tf���\�z<�Ah5X�=cL8�S�  
�Ai��>���O�R���e-�l�i��`  8!�Қ�ð��HfF� �`�RR�E=e�a��ԔbS�0Hv�� (�k��-�W�L*�{7�T�
37Z	<�a�k�{T��gmZ�|�=r�M��U[�u��\t�j NW���&�h����u;` �w������y���(|N�����bOg��`   p!)���A�����V:��%�C| 7F)��?�� �qZ	�Hh��3R�ĝ�E4aH~���>�AZ�n��R���r����`@L��Dǐ-���"H�$�<C�K�a��K��@.�u��an��!2� a��u��������6�� �  �!K�K�B<�.c�QÃE�Š�_(p��]Y� yL]�S� ��ht&ۗ4��R��c)r�>#0�Q�03,��c�eм1��ɇ�D�y����p4)�����i��/}�af3�g�6o,�#�&�]�ؕ���Zƌp`D���H&!���
�Ddۤ�פ/)iN\�  ��Zg�h   _�X��W�C���TP�9�W{;лH������bq�	��Hiu��v���tT?�����vsN
�=nb�Q ���l�6�w;��K��T�3�hζe���x����oy	��7D��)�M��H��i#�����8�F�-�W�[���T�A��+��v�pو����u����!�Q�����ڸE��s�+h�?�ۓ�H���<�*��S�e� �\J��Q�-�ț��.�LOJ�������`A��0w�ғ١�Pk�:��S��ʂ�#�o���M?x�Q�����?:`�T3�Hj�R��� ��4n``����Ҏ��V�%K�ћ�2��� �(�Q���;�8v�z �U +f��K��17�,`�<��6���	��.����Ph ��,!��r�W\7c�v���5������(�"��$�$���[���^����&pKo7���G�q���Iw������tә���6A<�y�'Z����?�%��R�OgC�@O�G`�Ofz�����+}�X�����K]��O����NE�,��
k���Ө�Gq��_�������GG�2�"����W�񄇺��j�_�_�t�F���­�N���G�:^�v�Y)l�8�Z�T��e�XYd�]��_ki�8!Q��b���~B��	�tݝPG+�P���@V�iw?��>`8F�g}2Wb멖H��ꃟ��� KmG^3#��J� 9��I�Q/:W`H>�6���Ԩ}���_�Gq��b�-Z�(�cܞQ�,?�c�}q��N�b�-��Yi�؟L
��lH,OI�]>o�ي��]��D��C~� 7��V��3�=�Q�	A&�3��c+�'N�/�%X��+�ց���T���8z�>���G߻Lp|�)F:@�-zx���Q�W�覾fn��*���O&�����¬0�j��Κ�U��K���A�v��J��=�����@��j��m(2̴K�ָ��䄥�#ی�#R*��`ʘb��x�b�8�,�M��:��n�IaY�X�Tn9�T���!k�{	!~��چ)[�$�>0C�����xK�:�ʲ��z�]�ˢM�.E2�?õ�����D�P��F���+�*}'�^+��Od3M�� ߨH�?J�Q� s�wH�dGn�I��G�W���ק����g��-O�Qޝbf��g�6�� {��	7]��?Bs��2�52������	���_�$��7B2U�;|��}�
�0�ɽ��p ?�!�׀�;�_�Ɛ{�+!�
:ǑYۂ� Ru9�UV���I�W�����XuT)ޥ�ŷXk~��>rWʅ�S-�p
̲�9�O_F�����3��2���?U2{o'��uO'�m,��������c̱��a;t�;r��x@4b��-��m������4m�]�G>u�Ҿ&�"�����v�M\�c�Rib��&�ֲ��y�iJ�WQvO9
�п�U/8��G��R��.8;8�:\;$=���a�e�<�vZ'm�脖+G����,\��e��&KW&l��"����2�B�y���e�J��+z/6euur�����?r$A�M6+nx)�/���]���O�m��y<+\O&��:,�3F�?���V[zC4�{��� pVk��������,��3��: 겾���u�#(��%k0>89���^��8�W�s�v,�x:���A���*��E7E�#|�ehuW�#���`Հ��a9l�{�������H�"��O��=�|�;껦5��P�w��������uK�����Fw;͎�"�E3Zξ,8�t��cf��ڤ��5�� ��9�k��~����k��+����E���d�yM/b�Ƞ����fE��	�;�Π�5�F{t\J�&�G_N�'�P�`j��«X>��dg���yD���4���˺��p��/�Tս]AN�T���>9I�k0]� �8��V��+MC���SIE�h�Іu�߶O��u-�W��E�V�@-��F���_V���e����䇕�/{R	OXc?��D;97�pH��y��}�s*���7����v�Eqr�d��>�\���\̵��#�IZְ��IUt��Az�!�g�xH�Oq�xX�W���&4�Ir��1|���f���Q�"KO�A!��S(x嚷Y�������ϒ��c�zm^`�E
�b��yB�n��p��I����;ئ
`$sUYu��S��|}>T�vLw��p,��r���t�X|5~��L���no@%���$��So�:�!ِ*Ș���`�(� �\��dmQ���W��Ւ��G�8"ٗ9� vd4&��F����F9���)==wK���D.��J�
{M�7�ashY���/ذ� ,�_ml��~�b�'}�рZ��e��GW0`��`Jt& C�8Ug֎�,��z���^�c�̒n_�EC�G
�V]���͖��+J&����61������$,T;��X���q�ʯg�	����5(��|i��m2��~��sd;�u^�����ί]����ga Z���;�����=�s�\<�YS�,)���K��e5�V�ܳ_�_Lf6w�^d��@J��V����C�[�4u�F�������S�����}��u'����y�z���y�N�}���*/��)��]	��E5��^�P��4�%s�Ϙ��~�kтH���Ea�s0����9����a)<��{8/M�}s|w�h/�n���z]w�t���lZ��r���e��J��wl�Rqv#��/�j��r����o�/���F&�Qo�w\Q7o��=:���Xe9V��fX�׌$�o�<��2ON@���PF�|��$l�j���$������$I��m �)-+XM�y�,��$K�Upқ�[���F�|ߌ�Z�t�kk&U���)G�4�S��4\��4)����ӽ����(,O��a��n��m�4�\��%�>�I� �JCK��@7�2ݸ��f����/��-����i'p�D��_�a�H�> G4�J�H�` �qޚ����ӟ��&�և�۬��f�Hx�C�H�5ޑ?l�{�F0i���q6���f����OX֓�
�j��M Fq��t1���*]�yW�Vh�T��%�&.�gm]7��w+�@�����j��K��E�l�4Y-i�2r�m����A�U$���I���y��Mw�j�L�oC*o�*�gW��� �+�oAvfb?���$�ωZ9�CZn���C-fKx�D*υU�R��M�DOc&|�EqVy��V�QB���� R�����i���"� R�~9	�����l���<B2�����^;�H�h=�B�L1aЯb�I���Ғ�&vCw��c)W��|���׶x�aq�������;g����5�U�C	�t#<z�_���u�BJ��x_J�������~فG�K�P����{5��)P�6��ȕkp�Xs�����[+�t�]5dqŰ���u.�}Y"p �����^%=D��D�h�i��ɳ�b�[	�� �ҙ2/�{2�f%F�_(7��|A�7#:§@����y$ p�ܙ��� ��	�\��ş)�A�,U0gn��rqe�A���?�d�S]���Q3�!b�&g8��$���y��Ι��h\��Xi�&�v�P�+e��ɕ��w�a��.����]��^�쁦}e$�)Σe�&r1�A���c ��2T0�]���3{dk�5�X�DIЈ���eFh`C���٨}LO����69FG՚��0�G��R�/�|񲽣��a*�H�6*b �{��y�f��UÍ=��n���h�[l7��d'��ķ��~�j<�t�׈��fb�j�lg
���A�Ւ�y�&g� ��H5Ǣ�����/&O^8S�J��?Iѱ=�w�,�l��ґ��!�8,|q��2�ğ��8G��niO����1�� �,3���ŗ4$�$k�$j�[kƴ�2�����嶢Ȁ�/�϶��*a'!��گ�Bf�O�N�W7)�G��тT��|c]��/`P�k�x��}Np9�		M�<��uy��ܛ�KD%�ZSn��֘��ӈ%}����+�2{�
�k����\o-��4�9���9����$C�����%�Z_�a��U<��W���	D7ڢV�P�,,?�r��SM�G\�m~�r;��t�ݍZƥ~i���a"b��C�d��\��y1��bDc���B��b�h�¬fK�i��|#�Ї��� j�B�����*C"�:%%v�z��>��2^�]��j_���e/���>��n����߹�����j����7�A���������a���@l_T6?#w*����P^���,�͵PV�ğ=�t���S�2'�ѯcW��R&\a����M0e�|�eU��]n	�����.B���C[#�?��QJ���ˠ�ux��`����7݉�	��aj��]��t(�#��e�_c��egPG��s�%+d��|jE܃q�t�]�O�4U�ش�_h
Ga4���>����N���W�ھA]������ ��*a�@s��J&��z����"YV��>}��u���\��P�	��q��G�kR\�r��L
���(������܌�������Y��V�Pߴz�;�MeȮ�z���(H�|����0tW�4#c��覵'�E�JU��,���s�5���+J��Z,��.08�k���m�����j�z'W&
�17qo[7�O/��)�ô0�	��^�G3�8��w:�� ���EA5e�Y�H�����J۲��M@N�?��^B���
�8�Q�I�3�h�f��f�D���k�:��(:����\��9�o��Y���e�A��i0{�5
Ʊ��NQn���I°�{?
Lb�B��������(�/�Qm�2'��_'ݵ��]т�q��*�8�;��	��4����a�KL��g}6�?2�n%f�"�j)��Ӄ^xܾ@�c!KX} RN1�0����ЛHL� ql�#bB$�=�N�����!����0�[����k�=���י+�p��<}c�:�ts�O�'�N�����4Dy��a��������? ���g�h9HQ��Z����,R;nc,*�AJ����UR#�X��_wO��nWH�� {;	��a�,2�K�Ҷn�k�vJ	/�ƣ�$'eeB��EW��I_�O��)G���W溹VR4�������Z���c��7�z2:�w���b���Y1�LW�AX�4�h�<\�	&Ka�:	��K�8����:�
� ���4V��U2�}u%��t�M3�%�I)W!	B��e��������KMC^v� }���=vw^۠+��6��+|����MWOi�ڱ��@�g�����t�v�s����ZOS������M���<��'�lJ=(Ԓם��F��Df%���,��rdש6�t��iY֣`���B0�>c��v���l(;#$[ͥ{��U1��m�����ml�,S�9�G�C�r&��������F	WsP��	���#�E	^�㚉S�Qɩf�~�+�9B�=K�X�rX�;��AE�[G���������	 U��`]��[�a����B�"E^ g����F���X�q��˳X�R%�=�v i̧e�4��#'|��y�P��)."`7/��"v��YC��"�:�E0���
��2P��{�6���h�E6弰|P��6�����*���x�U������	��G����T��q��]�n&��𝧀��g�����Hi��1�Dsٞ�S�z��C��B2j�9��N��%��E��,��~��)���/u��t|���y�VR��b&Yˁ�����O��a	pz�H/���,(���-�fn▹�SΉ2O�,���G��)&�m�@��.f��:��`ʀ�
�`kP X'p��l�	I���%ʍ��E�C��S˂�$]��SZ��\�Sr ��ۢ.F�#�A~>T�zC���$[��'4S�>���*[=L9��L0t0&�)�bX�M�K��E��5~4��<P���d�Iz\�d��?��BI�L�R�����o�ix�St�{�~�6���%���탤�����"���j@!
�"��2��zǸ-�X�t�?��$Q�O���w?�{,mU9a��6l��?|La"7��Jڀǂ��#�����'h0�ux\�	NOJڭc?�+�G`�f=ǝ���Q$ST�%�n�e+#L��Y/�FL��p�����MP��+笈�����~ڴ9�<�SBIL��f�P!��[����i
D�)M��`h����$��<HN&Q�#���(ػ��t�PI�JI��d��s7��"����I`+��e��/�q�!�˜��@�;4D%a�hS�=��J�&t6 ����⢛a��Hg�{�6�#��]��E��v����X�V"�����#�q�z�D2}��$�zLU�j�\���z���U��;��+�R�ĦwN���ơ����Ѩ�p��a�R�Eg5���]4�B�MĔ;��=��f~`7 ��2�P�[��8K@��s7�ԿKS�� ��w��EE"S��\1h�^�h�q��H�Pp`���"�O�1��5���c$������J��;d�e�TS&���.�j��i<?�97v���_8卵��Y�D�[�@�E)�  !�"'RW�c���ƅ�X�?
��(��?�}�Zi\_���r|��ٓ�>k��"FԶ]r��%k�����51�W|*��EN"�����܋��%�|c�ҕ��}���/���V��A�1�p�DDK+h�+D�|x��3E�i�����.d-$�@�{C'�� 'G����b��0M�3�ê��(sw�쾞����d������Y�bu��9�G\�0�	��2&�`�Ƃ5�/&�����+�0��P�.����+>�i ��4��bĄW�r!$�q0m��<��VA�����E�$q�];�ˏ�d~�q���Ox�g�n���\��4F�b�<A�&}<K��x�10���e 8��n�1l��;4u��r�Z��\�x�)f�e]�^�!n���r���uU��-����!�n����������YM�>攢1�w����q7]�d�7�@2���DEΣb��� 6͐�����Gw�i���4��.@A�)糴 �u}�ܭ�L�,�u���ڸV6�����
��`��k�@�J2P?����T4E�C��o�xy�
���r�5�@h�ZT��:o!�;��/��9��W��n��}������j
`��L�\�7��R�Zl�|r�m�x�Nr����H,�,�������7,cB_�����6�R�E�L�O��ؾ�8`�I��	�rE,�PY.M�f���+t +@aK�y Gc��*�lz���ta����^���U����j� �=a+�ML�t6ּa��I`A��?q�LN�C62TE7U_c%�¬��i��?��U׳�ő��G��p����nY8����G���ET��@�A(�6�%��6:���l9c=�7�=��A-1�4��L՘9���[��u�Q��`;�g���cϱ7�D�6?w�f"DfV��>��A�����3)]�d�\5��s;�5g/�h!Ӻ3��$���>6����<�O���oDĴg���M���#O<yN��;hz��h`����?�>S���N��Z	� �$���e�%�'d���~��j�r��=�bk��m��g��y"*�0Dީ��]�Rp���"�1�f>�Qc΍�ƧCT�W'�\�b J��{_�	dz����o/fbF�ۑ9K6��o`$�1w��>�����
;<�n���+'�B�!qIc��٨N�9���	vY�\�X�`.���Z?��	��$�łxͥq���Ĥ�:A�*C��⦽Λ��& �*��Ov�e����U��7	�?��Obp��2�@�ݡҍ�x�<KI9�D��2}�{}Zp�Dx�
�  p ���U�"��uߕx茙d���Vh�0��+lhk4r�Y��&9�~� �л���=`w�~��RH�*�]����;���
x!�����5��-�Kq$j�������e]�L\i��7	�O������*U�Tv!d_���xړe�����L�e�b�[&+R= �5HS���L�>
�b��{ԣ1��$�J�p�X�K�<�l��ע�/_J����(���!����
3Ā�I�[0}T���4�e��1��N������@3�72z�4�<�{z.��:� ��DV4�����NFLۀ�./�3���E[C�H�5i��Rj]��cOoH*y���ҕ���\[��9Ҡ!����k�O�&��Psg�����~�@ �b������_;���wu���&	fUn����l�{�Y�T.�ai�%�s��Cp�Q���èk���ؐ����M�����_�Ta+�D;�����B����"I0?��Pxg=��gY%��`Ue![���w#͎%5�&��#��	{:Y�eE�/���j��}:4u����i"z��Zxk����g拏J-?�(���hu�禜��36d1V󸁼4��}%V���BM�{��F}F�Y���1j� �1��GЦ��e�\��!g{��w8a��<5�r�q�Ƽ��{T���Ϊⵔm�e�?3
)2�$A�Jm�\ѯ�O�~r�@'u���/�*:,�J�(Zy8C�s�"S+�wo��*���6u��U9����y0qזW��/��|~��u�������q;�Ʌw�'�?&ou9����qzR��2��%a�NӲD�����R�䡃Q���CǼs�,��umM�љ:�jjSsO�?��C �������:�`�S Z8�Bkz������G����o.��l��6E�P7��BY�2O_&����#`pӏ��0��LZ _�X�� ��"�I����J�"W�q����d�JE����8�q�*�atw�d�g��^��� H�:B����5���P�/lCQ�댶�Ԇ(wB�25C	vp3R��!��V�uu�4L6���;H�5a�3�9���۫ؼ���6� �tqF��`֯TiT� �G�yUC�Cׁ
�   � ��u�!���є�he8�嬘�����@���9��y[�pV�8Z�ɻJ�z��}��Rk8���G�r]H�v��HE;3��#R��<U�L�S�Aɉ��W݆;wۍǱx���b��&�=��\ m|����s���fto9�d	vsԪ�œ�
��T����v��Y�o���^����L��^L1O����-� �$oQq$��`nH�.��|�&�{��򴨦�6�Fm �����d4`S��O��	;��˴6�G3I�>1�tɧvI�7]���{q���3��"4�]:O���X"��b�D�G+c��XJ��]�xu�/`;8��9v}�aܮ���s�|EpYc�Ve7�$Y��yR���hJ�6����N6��	���n�{Ic�rj������ � �BPNq�����V��L4���y��>[�A&�ua7�c�� ��w!v0�P���q�:4؅��s�zM�0������N��Ã+��/' ����}�ě=�4�l V���C���ّ��3L�V32o2���P�H�8h�Ç˫���$�Ȥ��1*�H���n�{i+`�J����`z�3b��Rs�G�� � -��Vd���I`n����p���W����U:α�7nɜ���I�E�M��4wg������)����P0��-��y��բ調:�� 0���ͽ<Y0�~I�]6�mRMo,:�`�)Vʿ٫3�gQJ � ja�zf��Z7�-����@V=�ںP)ռy9�^���4)H4�aݥ��\f��fU	�k�,���� a�[�4e�7DA0_���g��+w%e��:	CB�>��s[��Y���=��|�1��?Ú�K|�	ԉ�,0���z�N��;F���!�-��Hh�J�t���E�k3M��(��TE�O�z9#]���q�� �}mD/怎b�;�H��<P���lZPm�A�|x�A��>   � �B-���ÿ4��E�<�6��u��_�n5	c2��:GeDJ+m�j�z���(E���?X�,6�y��1R�(�}�'��._ť����W�1�3�A�\�[����F���\�/X�m^<	�<�r�NQ�#�.��Z	�m�4�/"�цT���=�	j�ܲ�K��a����
!�:5��3پ����y˶�̞���89����J-�(�S� �ZB^�(� ��$߳��$r�u�N�K�����*�T¤��1�=N`5�8�Eg:��S_��R�RtfC�l�/���<_�	�»"��O�o������%��%5�a������"�m��D��<���d��z��cn8H�w����l:�Sǐ�k���Y��*n�r�aПï��?5x��.���ߟR�G:�Ϩ�d'��Ռ��g#�ni��z{�l���1,��g�����-��3��K6���a!?�(�{,�i�C2���R�E<�	��������!y���± lLa{F �XVy4���_������B	|݋D��wC����YyfD W>'�y<-�R� R��/�cBX������(�ɏ�J�B ��?��~�� ��ƿ�SY�.q K���>V�/�$�e/������w������     !���C�hHQhc��MS0�E�5v?�]I��ֆ��
[���L��K�-,��g���LAǁ��U {��i�*NZ-��K� ��f�������_����
�ӓ�"�EH('�!H�"@[, �����x6�c���T�Sm�]��    !���C���(+2���PF��2�[��t<�\�s'�y[B)s�tA�L%��9>��)�`�M�L�b��)X�lUk>!��[Â�����q�HV�8��O,th���禦�'��pJ��(���0��¯n �A��!ju�h1��% ~3>���bPh1�8!�����&&����OF�z�5Հ�(c���m��|p1-��GAFI2�h#?��m�)�.�z�1ې�O��;�4(�y��s�Z�ͅ��?��+g��n�ܬ�����k� `?[�}�~}@KOdH%ؔYfU(��+)�^�u��Z  �!�ҚĤ��P"+
���  *��5�5e�H�T�]��%j��~������pl��<�kE$��)��ܜ�9����m4wy*�»ܜJ�-dZ�x�Yh��{6�*�[��P����`]p��N�Шj������w���V}p��z���  p!���Š�l!!B2��+��J���A ��{�m�y�ە�jir4�6K�I�Ϣ�ĝ:c���\z~;�$˷��7[DH��>ı	`�:#��a��Uv����R�3�;�JN76�T%�#E$���t�:6�F}�3�J�B�`8�U��:Q��!YIϬw&{~�h  !���'�XP3��#@�=���0;��	�*�~���+�w��Wg]� �K�K�oE$����`L�_�'�T��g\�T/1RY?6ơeX�C1��+�wx�2ԛg�1�m^���y{~`Uٴ{���&��=\_��+Z�1.�L�	�Ǿ�t�.C�X�X��:�i
�ZF���A�  p!��DX�1%��� U�l�}I7U�}?�Krd�5����3����� ��Ӣ�Kx��^�0���k+����|�Xށ����d
O%�W����~�ʉO+�`�ηu�ӠR��ס���:X	�`h� h~����)��P9������}q����     �V5�8   -Ѐ����C����l���G�x��l��Ð�~�VtNlN��	��)�'o���OpFg0��`�����[���9a��B!|_��ҽ�Uk[��Sw����*U����pL7c�qc�@��r��]C�L���,H�B�T���c��(*��lTZ��y�Rܟ���,�D�9.��/:b�A;��Ϭ��fߔ�:����l�a'&�(�a��RW��>���$��{���_s��Iz�%XQr��o��oNZ��&��?Jm����h��xm��� ��Ux5�����w����,g�ڢ�>�w�M��nd����X�?Й��Z1|�=��PYo)�\�wk:�$�d�M8��J#����}�Y��e�%���S#'��Ôuv��#=��,6#�+a��
}d�k�0�x��Y�\���dSD	e̕^����d�w�1�~�Ei0�3��J�#i�[�&8�<�0L���:����a���pG���<�e�����#fn�3]�}�����US�� �S���Y���%!A j����BS��=x�{kL��&0!I�^������Y -�Bo_��!�jY���)	��:��M�g+7��znNyP��׳HT�"J�W��%����0I���ݵ�b�\�����O�&֘��V�扔>�p�ҹ^%;7VL�s��cq0�-���1�_��(w։S�3�!�������gP�����f_/C8�1��,����{s��OOm��	;��b��YsF���b �YP���s@�-;�<��;�``Y�_�Ү��8�<��!t-Q�R��
��K}eM�D%�+�	L�C�y�_�&[R@J]��<Ѷ�ڿ5�^99z�����A '� o+�;@n��������;���2�.f;�������7��~޿-�թ�+W?�v%�+t]�>�7��G0��<q�H��>�@jn�1�l��Nd0�0z�=��N�f�A�}&yF�G%�X����O
\��ιc�־��$L�5�{(�����aZ��U���S�)p����qt�MdD��a���`��k3E7z*sfO�z�M�0��8�����ő7������%T�0P{oe,��z�J�D�+B�8�f�I>�G��Vs>r�L��J3j�-���~�2�?4����
��ܤ_媎;z?^�9R���h�?o~YHL��$���/^%��ݺP�(2�M��F���䦔��s(`�����;�i�v���;�hYm`�#�Ƀd"���H�?����bU;&��70	섚A����t]�J�^�M�q��F�,��>1����KԴ��o�vw�B?.�3���og�����s��1Hs,w��z�oj��c��������h�35�=W����,�p{�F��$z�P�%��f�y����Q��X�au#��5�)�����w=yN���X���o)/�"C�|��JQ,�b�u4Q?N�*Ɠe��`9-1��zH�3�Zv; �P�E�r��9��a���:�����6Y,���)�H�����%3���k�E�O�����PEq�'�q{������qѐ#�h��
} J+��~���{)�2���:K��ba��"��>�j�x�|��{A���z�8њ������?�m!�[�̢e���������ځ[�v����1	�6��8���n|���C8�� ������ܚ�(�v%�h�ې6������d<n��e�>rvW�H�N�R����O�2�Z���gGF��J�(I�	��x�5"���2��T}�K5�ȓS)�g���}Q5r�������S:��c�ڋ
��ҿ��.[(4� ]���6P��˝�V�<��fb�-�lnhf��O�q��NUG�9r��6i�T,y��.r�g�2�=Q\w���%Fy�ҥ+m�$�{k�s�2���T�$6������.q����Qg�1��K� >�З-��,�8~�����g.Y�|c� Ɩ�Z�7�k�=����O��hnu�"bg�ɹ=��!�A.�⩖��Ex������D��,B��t�Q�\0��ű�Ǎ�!~�2�g��h�|eDN.�:7�N�Uz���?�Y.���]���}���9 ����'6�g��p6�a�#����� Y�O�U��R"˛w�W���v���ZgڎdFn��oHdN� ���9Z�h����"﯁�x�ؿ:Q���*�G���D���P��V\]\y�Ñq��gU?�9%��- %�Ps��~Gm2��$���湭���%�S��Z2d�R5�x.���Ƶ@-o+޻��sK��U�������bE5��EV�!��Z2�=�E��		����H�tY6��x�mE�I�LM����j6x%��j� �O��	�+��"N�@�2ҟ�n�)��k�R�w���$,R��5�wI_�P\�F�p���	q1�/�@W��#_d�ZY��-!I ��8Z��+&�;Y'8�p7q����	1|	3�����4�-��oOF�n#N�dGl%��� ��M,��-���t����10(O].*�iA���;�p��y���-���G�G���%S��%͉����˾�A�1���>SR�t7Ɨ��h�&(�T��ی�����w�k�N�N-�6ڰ.�X�׼��C�M�k8���2"b�� ��Ò�P։�C3h<�͖ge� �k��5�y��{K�|�!�9�p�8�F�MoR��o~�c��Ȋ���u��ȋ��ŦOT��J)�����ytJ���j_���>��B*�pdi��|�ۃu#�q����)�LN�
�|vs�o�0Ic�h�K@�'�4��)�ݠȃt��SĤ�y!��eY���-^]�oH<�^9�ϙ����*V��1͛��9�&}C\sWdдG_��)S��ۃ��q����ʼ4�V�B4i�i����&�pd��S�*�=�s�~`_y����U�?��a+i�5=H�Y҇���� ��6Z ����g��g��h�V3�I?� ��q��"<�qv��� �e����3W�(������� �p:|@TY�a���&d�x���B��+�؁���.Ǩ��[����*M*,/^�iX�D�>J}rF�6vnG�Y���
�Ak�*���؃w���t!#�IL��$0�u۽"i!lP�YË[��-w5�d����@>Ӝ�nm���=t�_d����ג�}���lӑ:�v{�ň���wbi�^S=�
���m���8-�_��s��Sg����������H�5֣�T��5�6$��Jy�y�RM��: ��!�*�w��|������HY��N�@�>��Sy�ۣbj��[Fr�u�7x~T0S�7�Z�=���p$`M�r��H�����d�;�s�g�|�M�1U�M�|������E�B�:��N`q�h�]��H�NI�������h
�ў�\q�R�Z��=�'k;�O���s��vpG�:iX3{��UZ� q5x.?����G(�
�F�#�Z�����j���3�Ǔ.$c5M�#'��O'���{�)�r_{Tٯ��EUk���Q�cq
-4�exp��ɂ�������G���DP;��]dR��+�H,�uF��S�Qh���}�8���"o������A�u$�� [Z7٬����L���x�_,3�zV��/���>C��eM���q!���A)�k�dm��ݔ�Lg�-a�[J�٣
��tK��x��AT�H�>=�x��t̪�F�|0I�e�_�|��,���t�;����zϔ�A�T�l�59_����#����h��{Ta�{�&&sj��p�h��=��K�2�(Z����.�hJ{zK�q�L
�\XF��0�'�oV�jZ���L����_�4�H�r��}���X��j#�<3�ݑj�.�Q�X񻂜r
��sˀԆ�3!_ԙi���:iC��
����f
���/͋�����kb��!#~b��v�x��C��x#�7�jˋ�^�Wic;N�w���ǿ�E�}M�L�MOݭp/mY<��0Կ�CoX 9�B�k�%�G��\�
���C(����6�O�m��$��!�	,3��;A`JR𲮕�R}%!�f�Ҽ*E����~J�`18"���H9�U��&�/Uv������i�H�Ze����<��9�
<ҁ'ؕ3̑{~�_�h�C?�-�R3���P��e�LJ�|�ph���ݲ�S��9�H�CW��~�pY�
���#�ko��OɎT�1nM��t�E~�*��s�ڎ�dcj���m@�eT�S,�J������l�&�{�&�Q���}lf��\�WMS�x�1v�9�z^X��ny�0Bkxf`�N�gIEg~��5��Rt�ƶ����[,=��1�C0)�w��}���]�z#��lf�ը���"� ��Z/����33�z�.V��q��!,/�
 {�G�Oz�j�hu��CJ�J��: 5I��h����}���$�sd;��.A �� �?з(%X�����s�����f�yr�$���i�H1�x���o�0c��A���H�l�s�����$�If���2Ok�΀�G��{�K�u���>Э@q���n�B����^xa��K�$7�>av�M�'��l�L�� �ҏU56l�k���pXU��p��cj8J�(��d�U�>�������jDֆ��wA�eY���z"�Q���UY������r���S"�^�jYP�E���KΪ�_[���o)?���i�)7
+��oRs>: a�,q'�tUP�6U�������&�\GIYj.(�X�K�P\Ucz�J{�5�C)�dcx��t������{FI��Eo׋����k2���,5���	7ճa�	��L�����=�0�����2I+�!�NH��ѕ����:Ano��`�(�0� ����
��yP�����N}�y��S}�36_i��lq��Eo5��9
��?�<��[�C�C1���U�y%���Hk,��t�Wր�3-�mV�/����U���脏lq;y���v�x.����s��n����N	듪�̓�����s�j���:����S�![�ć?b,�x�x���01���eנ
��<4a����(�x�Cm��M<t3�xG�3x:�Q0�K��i�{�ɤ&N��@��5�O�j���_���̶�=
=NX�B���n!��g��N���$K෿��k�\��Z-Y4q�A��5�ѱV�B�V�;f�d/�Ng�_`?�߲8�\�����ߐz�)Ķ
����R(���UY�e{�0��9��Z�C�XPn�5����ʞ���Zvtu�K���gɖ��o�ㄋ�}�����o�f<u��f#_`�M
��SV�t܈�� ���L��� ��F���KA��?��Y�Zg�Ej\��ʖ���w5�9�b@��:�����x����ƺ��Q*����F/̅۪틅l��J\@Ab��sȧ���:��wV��"{<����S�>� H(�[�|a&!��\������0�H+ X(�u;w��0� �	t��>?���u��r��_����1N���Σۚ����&zk�!&��+a������쓏R�0��Z6͏@�Eh��  `��'R��c��Ri�y"/�D�G����Q�ri1&����>yI���>��tς��S���Ŀ�{����O��>8[���Y�۟5T������L-���֋�C�Y9Ss� ɍAQނ3%�r���xB+V���D�3���s�$^9jI	�m�q�{!c��{e��2�w:У8'�#,�˙�w��)�l���x��,\S�V�*K���#���'���p4~���+��A6�co-!2O����k�e¾�5!<0bX19H���|]�/q�m1J�c�=�u��Svؗ<�$�����@��D^H�q�8�.oZj�0��� {���bBG��_H��Ñ�z��^�F�Vi>�V
�+�֗;�y��5HO�I�]��]�tB2�
���f�Q�q��Lވ���l��2�:�vˋ`;G�����Ͻ���n>�ZL�BT�If��
N��+���G����AE��%��I`