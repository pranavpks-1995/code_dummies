��u#-���꺁(�/��Z���Шn`�s�ȇ���~�'�X���)��o/��¨��>�t���������	�%q�2�;c�U��mq���8c-J�?���-�f�t��vN����J���q1��j�G�W<i�B#XǪ畠 �@�d�����P���g|۷�>>F$�=�U�x8hf%�[��2�>]?�A)f%+����2���q}@�׭0��/��T����/e U��#�h��u�^���S�gy[٧�V������n0�Ј�؃�o����p.I �e�����CǇպ��ǧ|z���6�D�N[S&�Cd�S�pl��W�E��~�f�hW��FR2�'3�������j̭���]#�[�ʳ�����*�܅C NK�C�v�9&��Kp+X�w��J��Z �T&���V��:���s��ﲾ�������@blI5�l}�e�0�}���$pѧ���(~��hŶ�p׀�||>��'	*���_`��M^����ΰ�%��y��J?�I&�mQ�БFzW׏��d な�1�֘�z_�21�v����" �7�C��x�:"ו-�Ε�����i�=9�O2�����~��-_Ǔ:1���q<����UI�N�	"<�f��n�U"���s�4E��|a���,�Q:�-�[I����GKDK�S�q���s�Բ����}E˲���6��9Δՠ��c�_ 5�>�Q��2iGʙ�/z���ň�r�nO�a�V������[S~)C`��&j �S�O�*9|,��K�m��;()s��>�
09!0ML���Js:u~c,���.�2���f�k44�����A}����E3|�����_�|�?1o�W0<��\0(O����˰gK�li���b���?I� ��;\_ZJ�%�m���G��}�S�1�j��A2x<�k|ډh΀�V
�"%�ՏLu�?i1\Ï?�̂������}�P�p�wȑ�I����G��8<�FU�5X���� ���`^ğ}���i�,9���B�O��1��P��u�>'�T?���`\�68�����l�߱s�p���%QBm�_˺�T4T�QJ��
>��Y��g�L.2��
��i=�0�~�@4`6>���_�1	l5���Je1�i����� �W�|��/��	N�� ��M홷4�օ������G�I_t�K��)�Af�0d
�&� ��gE8�5H!�/ݲ�9��>9�ѻ���l
�G��s��QX�wC=��-S����M�#0��;s�lZfj������"�i�9.���n,�F�/���'�,�� h�o�pm��s��b�L��˅K�O�&$\�[C� ��[h�Қ����8<�I�K��ؒ�x�_�/�Fˑ}ZJ��N~V?{�-g���M0��k��r%(7���";t�|�(��=17&����K%��ض�eD�-u���'fZK�����۹�T�����^��[Y���[OR�����ȍH�m���z�u��o�ܡ~��)��X��gr�7�r���J��w�ۓ�u���?��%������Y$�L�l��x��!��Z��t��d.J��-ú����n�]3�C�Mԧ	�j����h�!�|G�
�!W@dMQ��`�X��#<���@2�ēc���ו��9o���$�DML�6�p��G� 8h@������%b�Q?������N��u��	,̞�ep�8�H��s��sNu�	�L�PtAf���TjT�S`������bQ�.�E!���D��-��21��$[�b9���dv��v�z�]3��oš��t�$���B̍��e��Q��0IǬ\�c���^�<�L�>��0D�	�4�9��/�	4p^x;�-9�B��u�%��N\�LHR���P�/5@Z�(K\��5�PZ/����%M�
vE��ϟ��b��XI��lU���̕���0
�&�en��'���R������ֱ>]6Xf΂������ ��E�&�58��`_�h�ND�tq�Q>�ՙ�5U�ϑ	|����uj�*�t�����7�AHX��0E�c3S@7�&����+��f���6��1�*�:�e](So-U=3Pق�h�Ԁ8�\&�A���U�0+8=��)���~�e9�����[\4��⏎��4.��`�9-rD��.����js��#�TՓ'l���1���4C��I���͏�B2�����&zi��ooVNw��ǉe�[�ǁ�e�n]Lj"Jp���V�c�{�����Ԛ�*����9V�y|���v&&чc��R~ܽ�_H�&"����n���U�6}��v	�i6��.m�!.Fktm;�LD��_t��e-'4-��ZY��j�FfȔg4��GjI1��u7R�[�v�-)}��D����jՎV������pE�Z| f���
�����F���_�5d���5x����������ӜX	5G?)-e��`{���<�eʝ�Ӹ]9NI6G�"�=���o3c
C�U�=�8�s3tV��Q���ۂ�߳}f�.J�R+�P �D
�j�Y�� i�-����B��ďH��:F�&����]�l*�چ�@��$�H�N���Q�8
p�L�N"�"���m� ��"������YB�f�,Ja,=YBnk1h�޼�¬�R"���1����=D������<S@�9�n��v4f!-�q�sCcqD��3�/�s~����ϡM*P�$=���¿��PY�T���r���~םZ����t7�t7*|w郿�bᗯ��M#�᝴�/��T-�0s�@T����h��t8��aT�z�:#֣����)�{�O)�Nz�d�d�����+J�-\'���3������̐%9[�CŁ�j&Kf������R#Y���a����s�?�8���p��O�N4)����L���]�;�4t�QI��*��%��K�߾YL�Iփ��m��4�V~ȶ��K=zp��Rs���EW =�
J-�MN�O��_�,<9�+Q[u�qH�Z���'��B	�>z�7�
Q;V;G�@��)p�\7;9�����#Y���8��"�wQ]�W�lH��2�3��%Ӣ$ ��j�_>�7-�w�hY���O���hB�S9�-�5M�>xp�W��l�7������]���J<+�t�1�N�#t��|o�ذ���!
��i;���g]�i�+'�Fʍ���}2�E1�7�6ϓ>��c^H�)�v
=nZI7b�uo�Z�~'�4�{/�%��+��#���WP)f�� `��~k�!q�Ⱦ�C���m4Zj�� �����~�ڒ�wZ��z�ԝ�Y�I��M�4p�S�ow�o�� c�}��X�66��U�P��r7�Ӑ�g�O�C!�1�~���T��ӆĜ1�y��	b�㌵�Ss�	�˸�c� ����^�o��:ċi��ۏ$_7��09:�*�J���'xj��ܼ�8kgi�,f��)!�!�F�G�,��?��li���q(�D�\�ب���1�Y����D�'�2�'���P`��Q�O=�PξWvS���z-��UߓF�׎�dF�����U����r3&�*;T��%����ۿe��W*K��/W �Z4T��4YD��C)��T��PzN��ý�Њ��ocj�{ĺ��v���9�q�X�(QXM�J�{�~2?��4Aǧ�<�u!��l���e�k���d�	h���X���:�*�U"��a��������F��c�}�-�~	N�=Y
'y�ٹ��o�י 0N�<�-��:/����L?DxŖ����c�gN�<l�qh�c��>^Y����Ě4�m-��[�m��_�:'���3Я�����|{Q8�^y�������E��4�˟e���+sv����dv��M�Swd]�T����фN֞٥�,�����(�;t�G�ŕ��W%���V�fO��|mL:���f�6��j�$������U�M����sd1�	�C\�DÂBCv�?(RZ &�sw-kJVC��ӈ"r�%�zG��r2�p݂�D�Fr^�U{�4#�K���\T-o�� �[1��:�	u�t)� :�3Э37yȸÅ[\L��j�X�5�Tkn����!��-�b$�]kt�T��N�k���V�]NT�Rd������ƭ菟$g��aW�x6eM,����t��<T�(���X��ui�g��g�)50����
Y}���W�=��,!�#��Z�Tn_r�'�`��"�N��x	�P��7�)i�42�#K�j�mL��`�d���&&:�JU�uA�a��N��9�H��	�����x�W!k*�_���cPR2C ���S�{�5�:7,U�b�z��G3I��I*wl@�)^�pÎ�$�k����	�緌P[���!J� ��g"�/9�X��dxHY�ř*r���?����V���$�S�@�)d��%ר)/�\2�X�͉���5�Ya76��<���C[h�J]��Eb�*��� �R�I�E� 2����iQr���n��[U������aȄ3��6a:��f�)�~�.�M��͈7����*zK�haUv�����g��u2F�I`E�ո����!��![�M:sP����S��^�_��x}O�
��'�^�aVnA�ꭕ��i(�_5Ba}3B��<f�h��&�Z����:�l��F�b��+�SZ�[5�V��D�� 
�pn"l��r�\}�,��2���b��_�<`L�f������r�}����wl� ���\�>�?,��Jͨ�i��:|�{���s�*��|?f����a�g.!�9>Ǟʞ�LkT�����&m% �SD�WY#k��R�d�Ъ/U���%��Z+Bν(� ����5%2�~��2��1�C�Ko�e9X �����WQ E�(kKE�L��ſ��0c0k���A��;��" )$�ڦt�A��`��^h'��ԕyN폨��@��g-�ҹ������M���W|1}zP��F��G4���%����[��e)�������ۥSL6}i���X��9J*�������g�9���p52�O�G�3�}���������q�u�*��%���i½ܶ����|	���&F�N  ^4V))P���hlb���k�w�Zgh�}H�.$�u�^��w��7��&���A��~��t�{�%�$�qҊ��n₱��N�]E���[n���$��#\���p�AdF`h��],?�����$2`�Jl�� Dm[��ZbU]+^E�m�Ộ�|��(YC�R� ���Ք t���B�l���^�n�곬�8���Υ���{WN.���J�f�bp'�4��@r��������ض̆h�?l��/���@#�7ϵ^�: �yE���_�B�ˮ�v�R�<m{w����p��V�p?�י�o#5�<+����y+��8��.X^a��Y��A�,�ŽD��H&5����3�0���'N�r���PM�9N�S��f���%F.�_�w'HWd�$����Wg��IH0��~��aM��b`Yû�oPKJH�q������j��8����_���`��homG험_{u� ������8�cI�j��{F��tS��FӨw������L�t����TQ���͋eM�P�CӀ�����E���wU�i��m��{��J�(`o�'7/����5_��ՙ���a�3�[�P�1�6ց�b�۰�R3Ͱ����S��G��|��B�Γ���l��q!��e�=��$iVF�K�{O�KdZ*0��?���L���ҿ.u!�쾝�!�K�r�Ǖ��xq��"8ȏ��Q��ǿ}9���I��MEq��q��J��,/��@�RfV���Ú����l��.-ŕ\T��=�c�Q��-r��D�E�S��P?K)��ڦ�˪)<)�79-Į~�p>T��5�;�U'�	�z�ڥy�#�W��H	��O��m��4�-�Te�H-�[e��+f&����_��?�ɕW���2�%Q��!�������fE��<��=����T�e��/�x�.�`���3G�֨\4ޟ��F4�nNY�փ�<�Fh	�ƙ��i���/-6�rӧ���u��u�`��'�}es��N��5P��)����#�׷"9�D���NP���f�f���$o�hV���8P�ך�+DO#%�_��]~y%����VۺB�.�V��gp�p�#9xI�8M��_���ǭ_��>@@8j����uƩ�۽��&��̩���RdW3��cg��ӻt�a�)���cC��cǐ$d�R�k-72k�������0Gw*ů��pc��1nnJ $x��vr���N4U�>�{�Q�E�	g�IwĚ60�{<9�9�__ՙ�b�E0d8���-r�wl\xbs��\3��x�{knC}�*=��Q"q��;�����]��a���nl���HH���?dT����tqr�)�t(��z�s���p�B�尸f�,14( �c�>A��k�ܱ쳾ڙ1�h}���S�f��V����7��k-;K��)�H�-�}K��@<�U�p�!�`���5���)Ԣjw�����ΗL�-��k�ޒ�͸����.��צ��PJ�z�|$�v~�'��e3���������{�����2��vN�±a�3��.m�Zk�[�W�I��f>����E�j�b�4���r1&%ƻ��v$�2`��A猘텁����Ʉ��6�T���o]��¨=L� �O���B�ٹ��hM�N�z���S���ж�)Q��42{��}�PB�)T��XQ��{���T�f�J�";|dƵ�vL$)�'0c�%>qDR�u���C4ᗀ�l�Ѕ	��Yc��ܼ��6K4f7����F%�u,�QT�up��y��G~g�o�d����|�{�J���̠�'HG�VzC�g~(���Kg�t3	i�"̂Mz���U[
�tJ��R4�P�6�=�4��|�w����H0�qkj�
T�;� h��ES4��)��|%�덑>�qr/	���CS5] .4= �$�Uݚ��ŽG5���5��|!�K�U��)�GrضO���\�8?F����B��'X�$6y焰��D_؝�s����;��x��Y�&�lttnЇ��sO
b��@�ߒ��_L�R{��)�<[��`P����Y-_�'q��vlJZI|+���X��\5��ΰ>����]Ҩ��,n$�p���wa���k�?q��p��^��i�X�E���|D�kNX�'O3e��j��#��ono,r^r�cZ>�"9������]ށc�J�-?��|�,`�h��2_/$G,��o֑\]�E#�F�K��!�}� ���� �h���={;�Nr�L�C�<�������	C]\ٮ�&�i�Wb�W*���3B�0^��-����x��J$XU䴦�W�`����Ѿi��2��
��!M�f���D��k��U�I�N�Ih�s�7n��� w��ڄa�ij��G����
���/K���,X�K�����z�C%C(��J7�n��DR�'*�S;���ɛ&���k���0�%tt��h�r�A왻���D��˕�@�n�Ք|���(��D:���Ѓ��u�������]��4Ş���2���<^`�R�<hob~�K���b���N�B+J�?��1@��}��R���"a����rco�E򶕃f�3&�����Nɡ�)*���g�Dv!�-�k����j��|���L~��!L����pO�'_ZN��I=��I�GP�8����ŋ��$=�{䄍+�
��7{{�!�|�2�b�\�9mX�VƆ��%f:+F�-	����8���,��V'D�,�s��L�8�#HjWn��79����z�.�B?=>�r]!�DG����;gnkW�p������o����L!�׃t��UA�l���1���h݌�S56"(+ ÑY%��e,������0t	�(�%B�k�a�/8MH��
)��&�xH~7 <��ɣ��L���K)�c�Kʈ��u�D���Z
GդV�t�[�K�0��/�U����|$g�����	�6W =+�����<ބ�
m]V�qO�'q�zxU1l!����!�H&(k¥�Y��i�a���'e���B�ϰ�]�I�����G�稵&��N�0{�WXU�	.����wl-�[ΜV��P�k�	U$�o� 0�l���V��2-Z�G��f�l`
�!��:��