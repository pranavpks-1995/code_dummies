��Ex[kt���Q@�AR�6   J �-W���$zD�&PĐ��i��j�n��)����8H�:�����h�i$��]���`��|����3�S�:^J�����mQ8����ά'��ω�_�+s[�<.y�z��ge>��@�G8�}u�c������^>�-�x%�ܮ=f�o��n�9��?���.xUx@z���p���S-1<�}��	+��Ks�p�\����3�:�c���=��k l�먲
!mR�NR��V!�����$L�cB���@�p7�Q�A}X���I��m��3��Eyody��X���$��b ;�M�f׃k�S�.��x�Ba,��i7�D��{�������!�:tRi@� 4��f���!�5G]ڝ��\��&��C]κe�,טGnL�#Mf0��0^*w�N�32_��<��w�iբ�'��%��eX�����8�Os��
"A��� � 
 ��?�xC�=ȄL�-k����o^?��\n�t��U�$@��    8!��<��"�J�  Ѐ@��Iɿ�/f:v]�^�4��'�s�ܖt��
�}
�n�����ETO�k�']P�c�#��A���l<���}�����GE�F	ډ�(�	�)� ��: u�i���5*tr�	c<}@^;B%�T @��aqUQ�)TkH@�*� @�!����D�� @nD�g�� �~=�{oN���^�SU�%r�U����*c���#��Z����jȅ}~�� mNR.�
:^(#�^	ءy���D��5�`�
����`�,��<�����.�� ,�5h���=#US*�    !����C0�Q
�(Xޕu`��X�;_�٣�K�a�pP�X;cs��69N9O��u�[~��E����BCVu��b!	�#n�)"b}��K ke��0�*4쐧H��.�ma�.�4�)X3~\�U�dG�}�%� �,F
 kr�5�.F�!MS�.���4 �!��!��&�Gt �
�4 q�A�-�d�$���zupŢj�2�k T՗1<>����#¯�)��S]�˨�~�#��}�=ӛ�h�a=�w�N��4�3w�J`6�<�9��`�P@$F
���[���p�pSo��T�Ñ\@`  �!��5%$Nk� �(� ,�ؘ"�#B�6��$�M&�m0�j�n1,Ԭ#��%��y�IY�1җ����7}q�J���[Q�B��u������������e�,(t���������� &O�B  j�a�����j�^��_�Ӽ\���yӤ�cc"�k�T�26$x   �!��<�&# �,��.X0`
���zUF�1Xk)�7ʅnA�j��+�z���ҏ)�<�m��d��fbRz�I��>i'�����;��.�o�J���#�t�L�i�$;.�b����bX�	A��B��>��ҙv\^�c�0Zd#�o�1UO:�-ô") 0   0 �L��1   �Ѱ��W�C��M��։�я
�k��n�UM;�=E��)g��������*{�?�n��:���?ָsmr{����T�X����Ђ��u�ۘͿ-.Es۔%}��<�A~���Z"H�פ|�a�h�#3���U{�T+4������� ��C[�