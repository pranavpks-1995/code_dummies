9z�,��E)���.�@yq����J�)\��!�0I��U�< /�Qi�#ܬ'��CˋoY����؇�`���ނ��5�Q!Y��)D(&L�J	�>��PU%@b(�# ���Jl}h�o���Igy*cߔ����%~B�㓻�M�� D<�� ��7
]��J�+s[{9��E�� �!��\Z?|�� 8�b���-Dϟϗ�o����AKF�ڬ��PK3 ���qM�af�e�?d�#H'��h�*-�+����sN�-FD��b`
{�7�5�cϡ⿣�v6�������a.��	\<P �s/VPcx^�����UD"��f"Qr���]Sa]H !�
X`+)X� q�禚����p����L୆qm�:�	�e�h���ƀTܠT,��5T�;A(mi��ZB ��W�QD�" �9�E@1	OPf�����zG����cѰ;�v�C����0H��%��_� ��4���ƨ�u��N��n	0 ��E��   ��В���0��3����v=�i��R��I.�H3��#'*�K���� �~dB��Eu4�W����݆�6�y���v�4	X�=E
��|�D�EL�s�*�b�8�l��<�1^�ߵ��0L�7X���@]9Z��!G�s�������2I��Ɣ�#������`g�4�1�~%�<��㫥@~�s�o@���SşT��y�3��a��9�ze�1ų��M���
�����eSb���3C�Ao�����ajH[������{1��\���h�F��6m��������n:��D0{>'��,Rh�s�,��n�|�4~�����2�c�o.������,�$��-���H]̳%ԤpG;^����,�2�	��0�R����-�>��ح5fѠA����9���[*�uW���ؑ����FkY\Bb�A�2*�D��b^�z�`Nz�EFG#��8�̋V�J�x^/ܬ�i,vl�Ўvu��,3�����5>~��u'~��?{��ؕS�kh��w[���k9<H��Eq�
�c�]��O��{��~F��
��9@U�X���)(���Kw�F��9�b��O�=S�-��3����B.w��ʵY|-�Pގ�$�HU�
U�oa���L��r�t*��&"r����:��v�Jq	�6X6��N��� �5U�RY�l�Y�BHX�26;z�Fq@��������߫��W�$%%0s�w��-����
��OU�&Ua�.��
�L�E�+#(�,vl�� �m���lIFI��g�1�1C��S˓��⬣eug׌�l^h�
t�C�!}��0j.gUs��*��g���ek��O���g�"d�94䉒�y(Xz�:n�m�2�+|�m
<��,�^Q�9�ʑʷ�� `h�P��<�?'b�U��ܬ��cԳi�Έ��v���х��w&�}�Gk1=Q�j�)��r�P�Q"B���8kQ�u�"<�_QU��1��oH���� �[��D������ %���m�t�`Q�J��K<)T|L$��k�5�t[ךCu����t��FJ9`!��J�Ky�&"��N�(�i�mr"�j�j뢢�A���`�֮�kV�P��i�x�a�����@}�鱯�NRW�;D�D��a3�0���Im_/��1!;Fg �[��H���I�����j7ג	M0�Q�o�=�k)?���6^��[���[�M�#ӪG2�z�14t�@a�\!���`o�V$��2��[�|M`��6vd�)�x?N�mUA6�M�8P�1�\�w!��������x�YTw�b�*��;��x�j\�x�(����o�@�n?�S���0�<�{/E;��,6{��*��Kc��8C9y6��%�#x��A� J󽾈4��<�J܆�_���������3A9t$xb�����+U[�df�c�^}�U���l���aX�
�U���݈Pf��!k�N���W:�?�V��y��n'�E������1ϐ�A|�N  t�'W_q��;���p���`�d�T!����W�c��R}���އ6���{`uJ�5e�y��~®���OΖj;E�H�J8��>A:�sp���p�sO��ڍ��
����2͠�[PA#�\fI��	�b�x��uc4�#��5��W$$%P�x���,8�
�}l
��'q?�;�-^1����r�[$IKR�A��EA���;@����ɹ� �qJ�~��]�v�����"�B@d���>�	R��g����*�WM��?fH��Y�`�e/|yyJhަϣt[%�3������hϏ-���fJ������h�d��X�����������o�5>d`���~����w�ߊ���:�Wh�P�ΣA� �   � ���U�o�0��AT��Q��2K�\��y����.M�C ������a!|�F�����(C��4��(�#%�e#N�&��Δ�,��̨�����|4(��9N�]�b��n�ۅѫ�J�"\��4�r��e� ���sk��S�8h�5�x���g�f��õCJg�x"T��?�ƣ
۾��P�]�^Z!�>�1j�?��'�a��Xy'쑧��4��׋��(#�e����h�� \ޥ%p�j��A�$    � ���u�m��H]!��C��-�@��U\w���wy����W���Ȩg�,�`����/������v�v����3��ʴ�O+�9}�\ws��_azkk`�%f)1�� �Gs�1���b+�?5iªL�]�|@m�f�^]��x�!����3��6��!�d
���2,������s�ɷ��m�}�f	����t�倾g�j*���K#G��7܆OMp���-�,u�Х|��*�w�*j@� ��PH8����{��@��x    � �"-�����VQ��4�� �ђ�`���'��/�jviQ��LD�
2�G��b�Δ|^�T�*��4J�c�/ӹߥ�l^��-�25B--���M�o�� �;?�:�^`�~%^r���A�~����Հ�oz�Q�Q�A

ӀG�L;L���A�h�@d��(�&��n>�WP`�Gl�r   d������C��@f���4��d~`�b�'�hc �	OA��Z���@U+'Ȣ����7]�"��U�N��a�ߪ���*G�؟���kɓ+uI�q���`3�|�n*d�:��\���Gl9(S����v��l�h�ʺo�M#oM���5�����t�A:��>�U����:��G�j_�Ȟ2/Q��B1�ř�T�����0{�	�d�q[]�f�~3��)x��9ډł
j:���[H5p/��{lW�-s	ƅ�d�Q����<"�^�Y��j�)ٟ��NES �L��a��
.��A�KK�9[�drbe����鿘.�MΥ�xW��:x��ĝ��M�JW*1�l3F@!�+t�}NL�@.���H_��\�)�GT@lۺCJ�-��Y]�*�ˀ2!mvA_L��|���.f�a
wC��rx������d��.�֊�f�n��IZ=Fx�GTǳN1�����P	i����D���;��+wx�����@�zKb�^ID�ؘ��tt�}�;թ��-5c�b��Ym�h,�Ě���@�^�(����0��y���������7NZ���3s`�~zk�ߩ@�k
a���<�� <��~Ĩ�9u�xl�O��͝����C\��P�ȬnUx꟣@\�=�^�Rv���z0Q�f��c0l�APƜߜBa��G�y^����K92���C1�k��D����D;��da�}/Xpž1�O����WM��N�&m�fvZ=I���󢹝�5���\�BNKs��*���G~6�����;��-J"]O�ȴ'����Ű��Y�:ѕ��\��i��Q�mk�ȼ��#n?��
<Dv>�ḩ00ˊɕ���y�UAg#S���f+�'#zo�(3`�/n�w�v,��|y�:�7E����@���e��v_�����`�b�j�z;'g�)��~����O6@}Tէk1M�[�;�RRoX6#+�u����p�OL����b5p~�/�T�d��s�k�(6�Ju�����;�PZHa�����'d��A��=֍���o�Y�;W��/<dz���oб��M*	4��ir�5H˽��ƨLy��=tu�|�1�d˝��}	l6���"e����l��ָ�FW�AW�X�1��)o7��/�vs�@1�J�_2�:�GM�_�G��Q)�r-R	d����2�g�J�8���ڄ�x�;R\�$py_��Cl��c]�k����]&yH	��=F�K�zh&�����~hΰ"��G�@^����HI�u�p*b������?ޭn1z�{P��<4i�����A�%�^oE�o�(��)��'�sy�<��7�<7���ۢ���U?��Z��tL��T�y���E�N.V������Ř��D��u�E�\��Su�G������<~��B��J��E!�/����O`�*��$:���	�����V?5�0`��D;k���{���0$��4L��PB�r�}���E�M>Þ��c�c1-��R��������K���U���9��j������	u�ESC�=(�	 �$���� %z�a�C�v,H�R
�+���go|�_0��q�Y]!:@�\P ���ܶ�ѵ���Wp�]����v�~�l(�Ac���ugR7�5N���Z���kW��Y%�����\�A�ϼ�T�'��t�$���8Y�+~=p&���ҏޝ���?X�]/���Wq�]2`�D���o�uD�Zr_78+��������	�n+VN��G���v���'�fPH�-�S-�=����c���$�l�zKt���$���\) T�`�Rr�oo�(�dp�>���8(C?�H��B�=/���y�0�(�rOv��q�"=��W��9BS��ƣA2�  *�'R��c��SC��*Hp�����ɵ0(j�7"�M$�;�H���r�x�$Ֆ��j������S[�a�)1d����Bs3�N�1����Z�x�ZyB���>P��mZ�{���B��e@	9D��.͘�,��˯���%� R�'�[)ח��L�!E(�0��$��Ne��]{����஽��
S��T�N�ܿ�|)Z5Ԧz�A�
��a*�ia��=���?��a1�p�.a�QI��\��7Є���'�=j"�A�^]UWt2q0�
��u��Y���bW��t"p�Q8�A��   �f�U�x#��"@�2�@�N�6����RV�Ĭ�K?í�;#m �fx�|޹"�;q���y w� H��\���'�v�i`G�g�6��	*FyC �Y6�Q
��Y�˞�xy����ąe�\���g� ����d@�&�m(G����5(gpN�$�-�,�z��A���L��B��̀oRخ4���Q�uG�B����2��C
K��C@r�]����������yHc��K�����(
 бy�˫�z��~1��{�̾�@��    � ��u�j�,�D��F�u+:J���i�����Nw$�A�"����lM�=�|��߅�@�����4&�y��N���z�@S)=���q8�_���+y��&�m�90|�k��`>Hܔ��F�I��9�\y*��;����L|l��x-G岶�
1�p��G�$�n���c���c��%��>cGT�c<�1L�?6@RH�V]vY����@�H    � ��-����8|J��FP��/���P�nUcǽ������d4�BMh �(s�����s�22Ԋj{����d)]��	0�FO�0��g}�jϦ>�����q�D�TzZ,��3�=�}3�p@���鬞qD�+���/r�o��a{��Ыʣ{��W�Π3����R �����$�����l�����P�a{)�@��3�z(
�U��D)�D�УD�����������!��@�-2�Յ���:�1�7�J1e�(��-8$��>n�fj�OЧ�E������F��۴�A�(r|�M��y�VقpЭ�]uJ M�X���%�>U���M���i6�y���������Ü�����4�q �A`��BRZ嵨,�C 8!��)1��� u��/�(#��Z��wg���N���`, �(�vc �3閺m�x�;�f������F��V}��9��� ��0JU*�� ���A
n���L.#]�pf�Iz��r>t%l� .��4JQH�.�6i�T�P*  p!�
8pJ� t)g���?�����[8xBhJ�}�e�M���O,�T'h���Va��rC�M�B\�D&%�u!�`	T̠��9���c�xR�Kqm�Ϋ|�L3��� I���/@VL�UT�\��2����}�� !���m��W4 t����(��w�l3�y��}��Da� OyR�I���w������U��<���ITvY[�U.�M7�`���u#<h (U�q0$D���;��|��.�a��1�d/q�<_�,�~��$A�1��w8�qtB���,{��0T �J�ٱ�_� !�1R1����ӑz��	�O�u�z�����He��8]N�j4��U��s��>\'W��O<E� �Y�� ���ˀ�H� 1c6�
{��e��v���}5wrc��\���;CjI���*���~�뻇$- ��j� !��)Z/��v��@�jh9�^����NZ&чdB�v�{�s��*�Y��v��'E���$s@�A:�8F�{�e�@e��F�+�"&A`	��B �&��Pj��C���@�>`Վ���}� 8�$n�[p�� �T���tm�ǉJqxQ @!��`\���eo+�e�(8y b���R|�O'T5�,4P)XE2K�Z