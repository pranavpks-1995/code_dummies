�O��3 {,��=���]m��%ܸ��u3ǹ;���Wڬ�� �
�}9
�K�T��_P'س�VP#�
-�!��S���>y}�Zk	�b'�����lW�Y�H�< 0��X��Ea'rVX��d޲�����(�ɡn|��7�6�n�����r��Y��|;�*��}��������fNy�������P��^�p�i2�i��	1��>�T�L/�,q�C>\�?���L��g���nws|̚6�DWX�2�R0vc�ঀ^v��#�&�Y�RB<̉	O��lm
���O��Y�+t
j���x��nޏ����7�BE&DL�����!���>�g���w�@B,�f�^}ŷ� �|���� �?�����; ��+z0�Q�bn[Cf����Hai,����|�/���C��= Y�f[_��a����H�,n����5��x�~�<ޯ�/�Ӧ��V螦�U��i�f�\`��H! 8J��}��^�nG�7�̦�e9�� ��a�D� >���R $FL�Q�gS�r"�:���2����P�j���܎À�:�3�2.5s��"�.h+z?�4m͸�$��>�;]��"�t�����Wq1W����x�L";fy�"�ŝ�."˭���z����:l�C��H|�ɧ  0�#��tA��h�g�l��3mvii�Q��?�Ύ��mg��.3�+�!֜�Dr��Qp�A�(��Kx�LK2:�����/۩+����p7�4��l�
1,N�h�u���Ns����9z+�4+��\	���8A(���x;ϝlQ1Q���RqA�����!�eT�'�;6A�,4:w�]a���|�2�����n�4�#�._d.gD��i�E�S}���>�+]� ���
Z�����̧J��$z3��Ⱦ
��dB5b��`�-�DQ�k���IIiҼT�]qtC���9��Nԙ�aQ�*�x��G�_��N+�߽[����G�cr�C�X��6����<��a�ֻx��C_	W�,�CG�C ����L�#�6�_.Q�k�R�����*��)\լ��쌒^��r�Hk�8)o3�Wv��1�ɮ�Z���#�Z孏�FKv�ǥ*�o���NI�_��@�-d��ru�.������q�ƍw��Ṹ�)]TO
5B��E�1�oM�Ro5��a�.9k p�i�5=����8�8�%.i �ҰГ�o�&�2&BGi��v:`�!��V�H��m@�ׄ������6z�ʱGP���`
0��[7��r��x�XC���L���kP&?�-�3zr94b����Ȱ������S�>���i�ׯ���=m��J��#����'�����m����g�nZ(��� ��'I�
X���A	���eQp(dԞ)1�.8�0g��/�Ŕs�����z�uA\i�"`���L�V���!����`��ت�7)���3���P6c�W�U���lJ��|���KT��I�r���Z��7�����F�/p���{���r�NU���C�oA��w�VY����B�7�3��r(�{J_ֿpbE�������վ<��:��q���RKe��FNw�Z��:��X��J����7���v����8�y������m�s�h ijo�4�b@&7D����Zj��=8�!��E��
IL~b����C����h��}!h��������Qs���f ��Yz�Ǚb��ĳ�\�\ۮS�E]gM���,�/V� ��h&
��E�  
 ���_H�тG�Z�S��m��q�ͯ8q����c6�W��Sd�R��U�M
��K�
L1��Z*/�8���^S(�����O���+agе� ��b�
�1߃bF�N��+���rf�I���\�:���'qf��;w��r���>fa�E���kYS���G���x���Z]��z�iV��)1���^R���޶� ��Ա�.�ݧ���4��DݽYX�'��٥_>��d҅�؃ʗWǁ�E�2[y:(�|6g�gv�2�I���I�֕����D�Ǘ�E~�4¸3(�8��Ś����)�C�pTb����� &�H�׋�������`-�oT^�#y��{�]OW%���>@� {�9"�j&���ťڨ�� K�c���m:�K�JN�Oj�&��x���;^]�Q �*k����������ٻc������TH����x*��!Ò�7��qv�#�}S�z�YU"���� �=�	��`e1���������