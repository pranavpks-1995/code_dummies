/�FB�E,�������
s���J���Aaզ��-
�؉[�&��;1��U�^3P�n��b�Dy=���BJ@�ˆ��~mL)�D�3�c��g�=����;�	�_�P?$Ap�	�?0n���[��=:��#T���߼�����n�s	l�82�jNFj��҃�\f�t�k�_f�`C�?M����PP(r_}4�D��<��P�M���Pb���V��Ƅt}��v��)�(�4�̺e��
z�&�ăA��A��S��J���N�Ǯ��W�u����B8'mݪ���S�ۭ�1�`�ZqVx�b�0�_<~��wϰ{�ڲ۳�n��������\'QDH�֭NOޥC���'	7o��g���7�G��]t�A�(+��.W�����"b�]������1���!M����+��U�`�8���z�u�
X�'��*���ڹ}%�)eB����g��:{#Ѐ�m�W}/�>IY)y�D*&E.�}rz9g F�!���1�B�+�D�oW�.�U��΀^Z��iIg=�OG��7���_{�,~��h��k0D�b���hy]�X��CT+�Ǌ��ް���(�U	%�f�������}�'SՖ��'G��a�^��K�u�`q��r����G�徭�ߩ��:��2�)�Hʉ��ڬ�������E�O�M�̳�6��m#�u��:�¢K5��&��F�=�U1�MD��[� ��Q�\\���������r0G�6��I�P�nAE�N�n��;��)�є��=�<�ҤO����2]�-uL#ތ��k4��$;?M�5ۤВ��wf�5�cK��Y�-#{��a7g����FƩ\�8��t3B�L�t��#3�7�}9�|禂��Zܖ�9����42��QU�h���g��y��ہ�ѫ���1���S�3�v�{Ao�VNb�7�enkv�y������ڦ#f������%�d����W�0K��aix �t����N�l-�/���}N���#Ox"e�I!+�)GV�f$�r���_��B�Hj�-LcQ�F�#��j�|}k�ܱ��F������oA'}���%`��È� %,oj$��c���4ϧ6��g��g�	򌍟� }3�~׃`���b2	��0����8�dW�x�F���j�נ�"I�� ����:��̄�C��l���+r�i�j�w�	�er�,���6�+�AƫѡC{D�ô@�B�cW�R]�퓫�J�xW��96��l�8?�cv�{�i�g��K�{���'N�/�~�~�H�s
n�6�>�V{-�S��ِ��!�����"	 �����J�e�ɨ���Ō�*���<��)鵟LX�҈I��O�2���4M��z���6i���Y���� >��Wa֩�rn:7%+�w���$ӆQ���� �}oC���g!���%�ܦ�V�D4�W�hV�~m��!���jh�z�4;۟C�S�J.�A�x95����)���,�@aH����D&b�6P(��Z|���'�mp����:~r���C���4�R��E�*�u�hҠ?�Ñ��¾��uo��3F*�:�,~K�����ѿlh���0�1����;���!>|�J���7�`�l]��4n��Čo%p|6F�;j��aw����L��UE@����>[��� ��o���c���T�������Vc��L?�$
��!&Ƞ{��p��λR�E*ѐ�o��h
fêQ�ryc�3���M�]k��zƨ�1����ݖ�D�qR)������N�+i� ��b=(��|j�|a�|<�4�l�g�V;��.���ZNjIa&�*�2��R`Q�/�z�q%5�,^���*:|~�V��E�$���җn2�2��n�4�eGiڼ��33�t�4��#�#��?������T�p/�"�h~��$�t�fK�J_�4 �v|u�����J��_@I-'���h��:��A��N�j����A���<K�@�EQ~��)T�al �PN퍭���:�"��o���J(��z�J��G�՘W�b�!B'�:E�$�n �G(H'���Z|�K�_�8�A��sI�^��c��l�B3ƻ$l�C�D��,{-�jN�U_�PӴ|�Fg���-�C$ A����(mwhw7<Q��c���BU��b�+J�H_Q�8��rp$�"�q{6��iq�Vb�Ǘ&}�:�B��@>�Bٰ3���dڅw�#]d;Tj]���[Fc�4U�)�V�> }մG�<?�;��=X���AZ4���Bw�#�s�K2Q�_̩{���8e�u��z���!�c�hҽZ*�3q���4�@Q-��ɐn�f`�LL��F��|� i�#��&߶]M�w	b���:�}2!�Fk��
@��|������QW�ʯ�5*�����-�G*h
�J3�T^�����5�S�a�n`�2�ń��U�Id�{ܚ���Ky%Ӟ��:��
KLݻ�j	*�+~L�����&APV��:�Sy7������t?��2vM�P��xK�[/KR԰�	nڦ�dX�� ϸ���b{�ǌO��Ta�e��5[ܦ�\<���49��$n�ꫂz[���)��C�K�a�a��}����H6��2����}��(�JxdH�th��Cn��57?,�<�f>rh�plx�%R��ry���ws�{Q��.2�#�E	���
��P��wzq�垪kj��y�S�\�k 4��VM�B���[-�t�PI��]�7��,�ݦ>������C�R��)@?� f?~5���l@��K���ѐR�E�$z�L�[ ��[^TbS�D��L�"&/��w�g�~���+Q�:���5�!�5�#�U&�ɘ����Ԅ�D{?�7�F?���>[N������b,�{v�;�~3��c����;����/��<@I�D�~��W)�e�I���v����!_���HM�I���A�MR>�Gn�o�-U�-�s��-��W����#��d������<CRr���yd��|pš��Z̔����e~�T�=��7{E*���-�%��y�����)l�Y��0��m{@�L��w[0¹dM ���5y� �Jv��3����;�� 2޲��O��Z�(�����>Hl{�:��������?g.9b	�E�L�F@ʹ��R����,D,.�}������dο��Cۚ�N��0���~���N���߻����AA����Yn(�X���HxUw����z��W��D �x�~��-�W���Dd,�L�n;�tG�A�������.��GR�$h��2�ZeF�͕�b|6�C&6����gl�%;�z/�@�������h��+L�>���`i�>M.W�!LFo���v����̈́��N]pjR�,v�(�yOUd>