package initial_Acquistion;
	module program (Empty);
	endmodule
endpackage