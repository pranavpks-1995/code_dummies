<�^�a��C�F�1���¹�4`�P��#���ub�C��#B!0�L'����S�n�RzAi~����9ǽ�Ȇ]>M~�Vޞ�!\\���?��k5�;X���{��2? H\��z�pMG�.x{W�m_�����z�xȅ����|�_5���n�_�^�9����t�M(��و>�:�ҳ���.x-j�#�����
՜vlW
2Q�G,(�(>�S:��v�`-�_�$ (B���PA��t�A�'�cf[��۔���!�����(��)��)�JD��� �a���E��G/!��I����7�O�,�]"�~�����	��ѿ�8]cA��/����:;���*Cj}P�ϕ=�B�l7�&v�`�E]��U;]�����*�<G������ح)��jo3�F��c.x��Մf }�:�L���5�Övm���D~ �a�T9�ůe�^Y�8c\q;u����@�uJ��_�[�o��U�1�Ӌ"7�L�u�y�WL����B�A����n��dbkd3A4��g�lb�ArNV"�[k4T fFL����)Pf��&�]��'�!�%�rŃy��Q��=�j����� �����?�M�u���y?d�V,	�_^LH6K�m>�H0����.x�����p��]�9�#�.�j�Z�o��U��N�$^H�9yLBd�j����ܟ3�~���(Љ�����J��9Uϒ0�fx�}@�m��ܗ�67�4�k�.����!'��MHӦ��zS�/�>7A�s���P8��]����n���`O��U����
��z|�ɤ�϶!^�����,Y�{BҐDuIzs�hC4RV�tc�(�����Û�%�bsސ�U�=�~ǓM�E_<�4K��D2�X��_N��8Lę>i���t�t5���G��ڄ�d$#��z�+
�c ��Kzb�
������_����gC%f�߸_]�́�w���4�d�m�e:k�4BI�~m��ȫ��YXN8k	�_��
�~���-�^]��Ư[�O�6���\��"R(��g ��4�f���E�&Sr�������_��߆Ӳ�p��4j׋M�R��X-f6x 9!���xk%�&���3�$-�[��m�{9Z��&��Rj	4H��E߂ �̻�����!��9��"�����Fi`X �e3�"F	����H�
`_�cS��&%���
�D6f�@�K!���{?k�u�>�˲����)3Ko�;$�٣%֍rv�k�ݛ��2�H��d�{��si^=�a���b���
T @� �����&s��g�2���	���ڔM�kT����~ $��i�ܱY�B��uLDց�!��5RFD%^XT.� :^��\���" �\��elg���u]���ë1_m�1ZU�l�,3�C�i" ;3�>|
4`0�iJ���&�ɩ[\kJOj�P�ZH$q��fL�,�� b �!��K߷�I��(�;�!� :k�v�y6Z�ɱ  7������A&���Ѐ    p!��= �"�T��� =����v>[���F7e�b�M�ؐ-c�o�m�
*����R�'Y��S�R�"�ķ�3\|��uV[��^HD�rX#2\%\<����$(H���Xʸ�a�í�j���^?o��1   ��u���t0w�6���-��-�=�B
�b(\
�ր�0!��5FA�d!-M�˖ � �j�|k��̹gt�l�ip���)$���U��4�VJ��A�0�E�K��P��#����p�����0��R��w��fwf%K��Yږ�u��ې�Q���6�K�9�Kꮟ@	&1� � kIWV �;������ !����
�������
�J6
`�6kY  p!����$��@ 7� �	�R�_�@�����'/��(���Ռ�g5�0����<�Vӆ�]T�TN��Y���b��Q���J����/Nݓ�2���4��w�PPk�V?m��Ɉ�8�?:s2|�T6)��$�@� �, ����Ժ4/_�h0wȻ���sսD 
y� �~ m7ȃHפ*�5��  �!��5IA�f � ��Ql%������WgJ\^Sw�.���b��7�m��(N|[�8�x�u��ڂ(�[�X�����*�]�h�v+�o��ӡg��Q�Ӹ�l)���kb��=�&���^��6�Ԣ&�_����K���A]� �CH?�!��ɧ-l¹�\%J=0Ґ�/�&���bVA��Q�H]RH,�A   !��90��""1���@� XT34g*�� 
������&��I�ʉs�A�q���\I<�ժ��2_���CT T�����ʬ^0�+�nx��0��B�� U��Z��%�	d@�!� �0
T ?Ӌ�n"�Љ�1 J:~?���� --x���o�1UJge*֥��� �   � �!��=�5���yU��R�s�cS:Muw���7��%�O52d) �x*x�4��ؖKHPH�z��/��:�[�bu�8�\�,�R�1��$ئ�#�"  XsV���m�s\�����B�O� @0ˍ���"��M� !J��2Ǒ�{�;�0�DA� �   9֑I�c�0'�((K�-�@�t�<D��)G(}%�
��}[F���7(��h[�pDs�\H�M�_��@�;�eu�۵a�n0���	Ax��j��L4�O�����a�uAu�� ����FY��,�ߢ%@�K�w�U��;�ߧI4b\?��q�P������W��/,BK]7�m���e��_AF���@��S�8Ė����2��uC��綌����rG3쏺���يo
�w���`]`�3ˌ;@F�їi��9���zDߝ���Zn�!2�<9��H�.�T�n���K���+�.4�Tc	�Z�9��#G7R?�c[�T���7�z�
�|�H�2�����5�T�F�I[	2�Pϻ���,:dH;WA��P��s9>y��!�iu/`tԜ���F�HX�waV�U'L�N����<=����譊s�[,��{K��Bl��1ݳ%�/Z�S@Y7��X���������,!�k%�~�~O�p�,����\�fd���*Ʃ�זKW�NN�ѿ�2����/�V4�@y�1o�_�^O�}��C�$��}`��SB� ��ȓ�������Q��Ōq�V`=�Ŝ2�R�f�>��2f�*�0~�DD]g��#��.;,������jǔ�=��mA����.�$�5�?&�A5ZE�KSE5T}�,;&�G�#j|i��95Ἱ!;H�>6؆��\���X��Y�ɢ�wS��.���Qӈ�bU�Һ�&j4<v�w$�67%���xN\�=s^�m��;lAH�ɒ�y���Fm[T}�,|Nn�^D�1��	X u���
a�~+ M����K��'��)�_"�<]}�c�;F��'Ay/��+#N�nx :S�����hp�iSBs�x�҂b�������������E�Y��2��� �v6�T�^
0l`�js*�!Ϧ�1�xV�T
P|[EA����o��H~%HF�ż���/��3{�1F�>���Kхzj��� �+�rƶj��hf������0�0��h�����#.�"3���v#�
֮#��8��QЖӎ�=�c�A� S  ��xc�����k���@�×�h3(�G7���;�J��~��d'<m9i���M<К��S0'��Őղ�{2ur�j��:��K�$/�f��@��ÿA�E>Q=e��z'��c���S9^c#˝�$��eX��@In��t�p��u�&\����W���Y堗_+}W�D�v�b��;���X�l���d"����@���V�<l�P��!�.P*hyR%�X;^�X7����E��W���pDFEaEn�")��Mɧ{0]e�ţ�L}���j@�@� *   � ���~�c�Hӈ&����D����Z�<5� 은��A���}� lQ�o/@Ӳ��nW1b�����5q��4�������e�N��v�?�o�z��:�Gʨ�I�u��t�]�/�hvO���G�Iqlj5�&�@�Dl�![�Qʊ�FB�/.X@<���-7�|����txWH�Ox7W�y �J#N�y@0X[˒���,L��a��iA�6D���@�� }    � �&��F:0��=ID �;��`'� �dّ\��3����.Th�p��%�@f�Cע���IMp�,%��z�8����7 ��WV�Q9�����ы��v�Ng:@�ͳ���CR�7��X[S���͂���-)X��3�ҀCm��pr���d�:<������ �����q޴L��EZ�r��������!��9�!
U�Q�i �`<��