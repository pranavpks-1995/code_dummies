@��ڏv�޷�Nؒ���㙀p8��LQ/Fy�I�i{��6�.�R.-tۆm	�*8�)�{��u���5�wh�B��9tz�ҿ["���~���F�-Y���(sU%�Wl��)�"�@+Z��
G$/d�p�̀QU�`��3�����*)�����'���cY�ldZ���D7!�B0׫����1��!�2�Pu�� �]�b��w�:K��V�1�0�ZKC:�%Ӊ�0�_����Ү)3��`�pC����L��Uv7`s?0`I�v��k��%G��U	u�!�A�����yF��� $m��y�}�aad���3���Y�1V*��! ���#�cs�9���Un!����	�]�vS�9��S����3�;{�����I�4��o7s,ɤNs�H���L�?��nnk�L(^=�I_=I�6��SD��&�R���!*ҕ__f-������@+��n,r�B(���l����-��y}uz��)<Nent}�@cn�C`��PF+h
ϏyU���a����|ӗM9�Z����d��>��;:o��q��T/R>�����Hf1#!S+�b�ZYl})d�9%�i'�x�䡲A�	�܄�>P+�r�;�kB�?z�"��J��m��<G����*Lm�m*�F��hf��B��6Y��K2��$p�3�P�q*߾�j��B���>#c,�dH��+w��sf>|+]PzFQ�d���PA���O#Z�j�H�3��&R7��T��-*[!�;����s���M{�|�Qj�4�1���m�4�b^�L�Q��H�D,�  $ �����,t`��DV��sG����iN�ݢ��M,�j�ʢ�������=U�Hں�Hİ�r=0�Փ����1c��E0�r��*��	���T�ͼY���#��:�
�:���|�3�8�P�C���2�Z-dŭ�9�T��!��8���d�lx���Y�X�8K�����,ٌ�%j2�����{N�Pa*��qs�[Ȓ�#Jo�]H��\��,�M�K��^����������?B�d���r�V1��@��ԟ���ɘ��l����O̖�]�����2�: g�xxL�@�C԰q�DFg�6V䂕z	���\oΕ�Wh	�+���{1mZ6,o�^KU3�(���/6������d���H�bMxN4�������y�'1o����:a���^�i������O�q��W���O��5��^��]:F����[noD@���+G� -��3���z�C��r%|�|I�f�ĩ�q��
2T�F�y[ѡ�wY|��e+�S�z�����cy���y�*m�@����yS�|y~(�ҫ/@R�2�R�������$L�%KB�}�0SFj��m$�X8Cf�,�\����2�?>���/��ÑZ0��مRU+�#��>�n	��ȕ�u��R��O�u�Ż�#�|�'�H���Ja�q#��tU��Z���h��L�e�l��������C�ޏ)�~eY�wD	L�����g�>ƀ9��Lo}�Z���L˔�F �Jn��:4�|��-��y���m/4�c�qt�6�i��w��1;�W�y@p��4���_r������ƹu��}"��l98��(F��S�5P�g���eb�1�N	 � J�s\�}��6�,�jr��{$/5�)P]Ɣ�8��,�T�����p��l��W!�
�����ynk��z�9� �L���M��zy�>a�͛��|�l����������1I�{�۞�Z���
W3X+����qtƈPԂ�q+R���n��Dʹ�Z4�����U~@6����� Dm��EΦ�qè�H�I����AZK���9�����/g�m@�[�D(�a     �-W����l+K�jg�qpI�����	OpV����R�L2�C�������h�E�̝{�9���4y��޽Í(@�l�W� b�@��� v��J�,4�?i��������w���䫘�6���l��3aK���;��^��Y0��Fȼ�"",:p%K0���2Ĭ1<Zk��X,M�U�%�j��hb8���K$��Kt%5\�^U���f��������Z;S��l��ץ�&tIo�������e�
�8���M(�1N���� ftge�{���!��R����'��L|gֶeF��8\��h��0��@]���#b(rOlLo�!*p�|��\&M�����k����
�]_o��8=�+#��LJ"����L��\�L:Pv�F��
M��ꄌ�ѻJ�����ys�'$����hh�ۤ�-E�?3�.T#�"Z����=�v� � ���3]�ʈ��{����>"�:vb4x�u#�L����T��~C���`�������e��S9Bq�q9�F%�tj�F%𥽗��� �Z\�}�)��:���Bl�J���3���ajQ����	e�vඒ#A@��"3�Ҩb>r�����Ohi�u�]�Վ�0�1k������V-F1�FK#"� 7 ���ǅ�)$�t�F@P�����2$&���G9��x���ψn�V�x�D�,�K~,�>)��9���\��{����I[f_���^��Ч.!ཡ<<O	��G���4��!8L�H)La��M�+L �8"����;o�p;A�~���TMo�>�x 5z�Ul�H�����;E�mcXDT�hH6`����F:��W��S.8��t��~��>#֯���<Ċf\(����*�(Ղ�����|my@	7$��x�w�p��D!����G�'z2�Qˡ�=�%u�1C��ŵB�t��
�_$���T5��6�3�:�8m^&[aT�`��?���5N4�:�o�ȲО���!��KI���s@��s*���t�Z���q���C��ix���g��Ó5�j@�r����9U�H �EX���������!�������T� 2L4ƴ[Vt �ze�}�l10�~F���:�8���w��+.+�Z�@ E�G�<�� _m���b��o�ݳXWR��c�n�CIMfx��mI�zV�hno���.Մ�0��	�|�� ����o�?uQZS%�u�     �!��Ι��uw��k��(�ݲ�u��եl�s�ή��rk����?�ͷX;���6�4���R+B>��.�Q�ۖYTU�����ݯ�>M��H��g"���3�ZC(����Xӛ���ҝ�v-	me�j�Ծ��S�^�������.b�A�|����%@o�3uM��Y�P�� �    �!���Ga�Ql#
��ڲ��V� -A���CIZ뻚I��B�B�i��gɰ��b[d�s.�D�a����;����Vac���/������e��U!��	"������3�f	˗�z���e_���y���kd� �t�&D7yg	W�����	�\D

w?LD|6i*\P��T  �p!��@Z���Cv�Z0^�Z�}���pKh؄�٣�;�ld�3(�	l�8z<B����I�]f�냠d�1����f*�f��.b��y��S*ww�]c��1��F������C���ߺDu���M��xZ���ɒwl����p1O�V�}*�*����N�{,ϐ    !��V�5!D �ՄB�� ��ҭw���BB�q��������瘁��F��sU &�w��kpf�\�����з2)|�k��GG{�4�6��Bܒ�p�`RGx+�bXak�d�|(i0SAN�\h(�_���"ƫ�{�4�rA/�U=w�i}�_R��%N       8!���#� �**��g"�@$)E C� �����}O�.�)�FA5��R��c��۰҃h��_���{�Mr>����jD�x�7��ʸ�OO���3��7
PkV*���r�!�OQ����n׽�:�>G\�Z$�JS�����K/T��R����   �!���lJ+

�%"��0+9hJ�\j�,zO<�!��5ڐ��=�J�� j 0vGs �WPSK�Y(�y`XVK�n��֔�԰"&W����(S�4��%��Kv��O�8p�7�.m�7�	,̞:��
��B���eB
 �8�٫�/�� c��&�-!	L����ϙ� �!��*Ă�l��f�2��pP I���9/?�A����L�'"��H�����J�:'&nѪ�	#���>O���XŅ���g#��l�v��+>�(7d���d/n0��N���
Ž�@�j�QHXN &P�D<�|����ʛ1�'=@  p�P�1   �(�UW�C�����u�o&oC��=��N������ ���}0��V�r�m���S�(��fݾs]�����y����Wyވo�4ݞ9�9�C?�����)
\V]�Z=�J���;�;�V����P@��Ebs��덭J�V�V�?����+��L.ܘ>r��>����:��?9�k����y���On��A6�k���m;^���S�QW�K~ˉG-�ÃP�b;�x#2#4��/����q��A����H�]{B�~���lpGD�tՏ��χ5����c�:�TP�Y$?��N�r`��m���n�/=�g�2���b���2�Օ�2�Ӵ��y����jYМ��O�UV��e�Q�X6�j_�8zֹs̓�Xhv����>@5MY�y|	��3��";Ԯ
���<��s;������x���z���<q�4tf�?��2�J�W��mR��R���aףRD����R�?L&���I��8@�rRGxF��CR�UO'�<N�%��+�V��z�'��I�.0��C,�Υ�xV���xj���T�Ș�C�M�.y��ڏ�N���H��6k{?���D4`mt�����y��x#F4)�SU�Gx�G����}���N�!Q4����Ck%}�hK��h�\�c��Z]�ijD #i�F>5$ ~<�!C=�<����HOȫ�b�ь�,�j�ۈ�h��(�)3�6�4F3���9���h>����O�%���AU>Z�l�����LM"	 ����TAʏ���m��9K�����R��`�~g`/���;ǎ��5AB��]�Ha�ѐ>A����e��q�ڀ���!5V1	Qlۃ�g&^�� �N��O�a]z$������:���77�v3:J�
�*�Dt��Ic�<�䄚������U|��!"�46%8�4e�B^H���Ot.V�!]:wy@o_�Q�=�å�v	���?F~I��8���g[qE$�������ӏ����ϼېuI�Ð6U����~�?��ࡈ^�s�rP9M����p�/��US�-���^�Q� �Ϥ�z2�Z�C�%dZ��u�B�W~#���8D�1)�QXq2�eJ???~m[ ؏(���Ⱥv8n����Ǽ�y�H�h6���F��\�8�,�fh	�'��?s�eiM���7��(�c#��r�����	��~d�d�%R�MI�� M�ءd���_���$�Zd��� F-Y����܉�R����#�ΝZ�������U�ﵪq���}Y�ä����G��
�Q��3#!˿@h��<�>�s���/Q��8զ�=8�ӟ
	�Ѡ��Yf̛<�ax�p2��;��P�	��{:G\J�� (�uǢ�E���h��TV�Ɖ������9���gx�˴%13���#��D�(3r�u �9g�_�by��oe�p�\$�A�:���:Q�lg�+ma~�S� aVTϒqZ�b���Tb=ʬ�2`?b���/�\}�p����fL���*���,�؀|-��2פ5�S]���8�ŗ�Z���[�]�%9�au����H�T���u��B��/�
\�>\��N�	[����#�Pz}��'���?Nsf��rV3��<"R�h���ܮ���ǚ�����-s��¸#Ѥ&��Y���8`̷�+��#&��~ �	��k����(e�+�6e�O6H�����i�z&�5ݯʮ�2Ѝ��r>y���f�o׃��̙@�z�Qy�C�H�����"�nM�ve~_�-���Ȉ����o�d���\s����[jm�$�ۉ�8#�[��O��(0C��*��[��},R���$�\��NZ�٦��A<�E�2�DQ��b�^\�7~��.���X��l�}��d�)�p[mX�ޗ����ϕM�DhD�s�@�!��!�������R�4&�� ����<��=�l�͇�V�08���Ude9r �,i1Eqt�x�b"�n��tB���w�m P�=��Wq��
#s�t����)}Tʼ�����4�4H}��xYB��������N�X r�{�I�F�9�G�̽�ϓ�j�\��{nW-i���z�yEno�%3'uS8��$�����?�ȳu���'y�G�@;|�`�Lb�}U9C�1��P�h���Ͳ��|��3�%��Q�^�t �J�ST�+<�x���!��_��۔T�g�v��l���x�<󚡉��uĞwfc�4-����O�)ka�Ur'O]�m��Y����
po��t�H��Fw>��c�����瑍l����9Qhm�w�)�pж��~������̢����_0ZU�8��^Q���5��M�g�n�4lU78����@0"�2 S?��Md�W��y�Nwlú��	L;L�c��7
�de/U���W�&�I3"a*ɪ~B��K����X����_��>j(eiɀ�ʆ�	ԟNgj�SM#J�ܥ[v~��?̋�mTOg|�`r��۲"���)�0�7���	��AZl�l+�Z��c�����w%C�u��N�KD����j��%��%�#d�G�q�!�٘��^� �~)����Q2A�à#�+dԵ��37���-��C��3�%n�Ao�s{�W��L��}�_�'�zk��<U���#�Plh��r�X��tU�d��Q,�>@'rmm� �+���ۘ�W,�<7M�\�W�'~�u�|��)ρ�ٹ[6C�Ru��;~u��0��
��q�M�8<�&��+��u�ߌ�mWb4XAzF��H:c|֎�BF��(2�:�`��.���
 !�9�Y*	/��0�8�>P��0!�mT��	����&�]U�E��4�4�7�PS�*ƀ�jVI8k�1�\Y�:�<s����U@��:�]#�g�l~����*�2���U���m�x��|����`V��s!귫������FUo��~(ڬC��<~��� Џ^��3�^��$�^�:�d�������5@F&s�	�z���(�]�O\KJg9���l8��VF�w�q~q�k�p$�ki��s�c_򁈾�O1�݅�5�7���r����C��~���p��%P��nժ�N�A2��2�5��Ξ�ŎxD�/�`�|쯽^�n&
֞0E|�j|;�g�P���ᛣ�ń��5�l�$PR4 ص�<�p��hAˉ?�h������#��P�/�"�Vְe�R���b��Cڪ)��}<2t�,��w��́([�qy3|=�Q/zP�����S��"��G�|�$%N,B��oЙ,���ݲ�@�����ߜ$�-h����l�uö�l">���Ec�+�cn���XH2
��{8Z8�B�k��B��S�A4=�;WK}!)���&�,�SH����ۉhq�S�\���bŰdJYt"��OB�~�ܗ����h�ү�3�`Ϋ�ݹ���l����S�ZrA�'��0����^�k5	!�0��p'Xf'I�C�ۿo�F�'� 5*8G��W���Z�(�G�v�_���nN)���Ɔ��*�Ŀ֨��v;�}FOi�js	�B�>��/6�<���"�������	+rd��U
��m�|�L,�b�LF���#��ޓ'��1��:�\�*��M��[��T&��zQ/��������iv�q�1�0Q��d!XlA�2�P�'����#{�<���z�:��Nw��� ���o��.2�\����׀��"��֙w�u�p���lH�3ţ5C�oS���Ğ�b���h�,�L�-)�ԣ�#&!̵����n��BiE֨q�֘��[��ф��:�{Z�;GA�@�T���1��'��͈��%�Հ��t��?��$��V�}����?�g9����%=dէQ�#�^��3����,�>�D�Ŗ�Y����~��ha*q_t��r��C���x;ǯ�l�+�
)�M05�[rF؆FI��Z��6O����Y����m]��VM�Ϩx�^�������?Ƀ�Ge�R���5e�Mǥ��@��+�����5����6��
ʀ��T����O>d�GT��  L�b%RW�c�����2���&���=T��I����:-TR <��M�A��q�[���_@M׽��R�=�?
s��hde���:�^+���W��&�N�'��{-�� ����F/U�Kz���R~�^�\T��uM�mI��� ��8�C�Ci@��)�w ��Y�C �s���-���F�v�Y�%

�ǵ�����쨬�GcL�n�W{��[��b�$�Gty��x3DD�]2�-m%�!0���ݽ�#�&�I#�n����iÊ�G��ʒ�ڀ�G[-��-ra������D���
b\�~vP2�~l6���85�izG�/I�l��m��T�"��Æ"�p.<��iO���٢�V����5W�A��:���l�)� +T���U�FLrYg1l(��#U�mD�gIY ��f��D0F�������V@B�sN��gH�,�}!�����E�A�8��o�lI%4H�E���q��3 `�yQU|���۞ּ;OУ���Y�|{���-��.�g3(��F��0d�Uo�>��d���e�il-d77r��<ƺ�a�$L�Cat�g!�$��v�(�"?^�*�js0��"����X泶��ا@`�R�Z��8�P���w��%G��ME2ٲ
q�d)�y��� H�Ya!v5��e`��3>�7��g�J����d�i]�Wi����D1���4hS߫^��&^���c$�����'�*TO�~���}K�5� S-���:���N'(��,E\�Z7\�~�X��KJI2e�e���;:$�2�kR?ӗ=؅�S��Y�C)����V6��9�1�gO���e ���B�*�u���u�Wu$�.� �sa��i g�1;����4��ў<l����=�ɜ���<Z��#+� �;E�++�)}�"Lt�tˤ�x|�l�V���V*_�S�H�����G�lDeZAнe��Vԃ���A^��
�� _嶾<� ��k��=�,u��7���l�l�@�l3[_�y� �v�W#�Ϟ�:ǟ��а�_��J0;8���+��Q���u��J:a�B��GRG-v�nTL��}t�,�rI:��+����*Ƥ�.c�f�⨑�)+<g� ��%��~~���{3����������@K׿�󱼷�5{ߕ�K"��X�2�"�:�2�p�����X�ˋL�K����ռ��bs���"BO���E�Ww�����"=�R6�W��mckm���T	h��S�	M�K�[���]NB�5U|��R5�a�7�d�V���ٗy���h�֨�;qFQ�^���z�W���.�ͺ����}l��!)D�)�њ�z�^�
�j��y�����B�������/�����P �OF_ �j�J�q�8ڲ���j��ܟe���9%���i�Os5x��#���Qn�X2q񷙔�i�Z��<.�v���d�~܄����"n���Ӈ���w,�@:uu�y4f���A���bɂI~h��6$����P��J�\�a7�-T��x�"�+i����FM�l	�3Y��^β���%Y@�d�3O�:qS�j���H��W�aaY�7&jWB�)G�k� >�qX����ͥ^HJ�����E��hN/�͌HD��V2���5�-�q�V��
l�ь&��aX(<�I��w�RĘ0O|�&F�NW���Be��V��&o�_R=�4�M��iY��䄫L
�8W���5��3�\��`ߨ�(�*{E[�Nt@�wph���릘���zW3N��ZP`�2�	����zXN@D;B��D@e��:$��ZJ�l}����w�_S�i�oׄ�^��t���Q�����W��Cҁ�  � �F���,t`�c�GU����E����
S"�
��>��������$���\w����G�����W>�P�����a�¸�G����|[��c귾�Ε~|�yu�>��F��F���\�2h������'�/*��hB��87h� �Ω
���}D������V�1��!�fnv�$|��&��ϑ�8a�9�� P��WNw1��m���Z	�ҫ��Ly��+~j���0�F���V֫k�^����z<�IR���]���{R
M1���s#}��ːæ���3�D.��{q����V�S�g>Y���������>���e̛j�p_��)�U�r6�H��L)-L1F�����9��gz5:�sv��NY@�:ݻ��Aj����?��|>�h%��+��Sx�MY�`¢��OL�1%��+�h�ѣ'ư9�zS<*��7T����� ���^�T(�`�_��zD\�z�{�����ğ���i�:9	���{�ѾE����%V�r���;���i�*���!8b����Xи�����'�G���U��V)�3�ؐ�(|� �x^��ե�OD��O��f[$,��]pԥ���ϯt�Ȭ�_<NC��y�L�P�D�=C�����i�SJ