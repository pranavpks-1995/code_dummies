
?�&ɮ�~<Ti��w��ΟdF;�w�jF���tv^��N�5��d@L�q���.�Ü�Mwĳf�|�a�N�*��7rG��q���'�wn���Qn�S�*��d���<׾�Q�����Ix�8��_��QX��`lR�SHո�UEo��4�j(YD51�\6��b�`�e{�3\M�6�JXSB����%b*AA�R�/ᳬ{$$b���JPc��D��6����q��P/2�.I\P�8 �~����g��:�Jc�HB��]�o��N��#�}����6A^�6ʼ������,�Ǹu��|���^(�?��f�uk�AkFT���a]�(1�Z�w=�a?r�h��.Ƥ�e;��+�F�+��XЄ8�ZZ���E�pD�ɂ��p͍��4���_ȷA�l��s@12���o�i#|�ڙQ���Oq<)�S�@�z0/Z���ˎhC2�C�5% D9����X$ q�Z�1�)�J�y"ˌT<�
�D� q��4;�\Z�B_����*�X�t����xWS���=�;w��v����V���ݤ��Pc���*���'�{�G)�I �k���d� ����P=-��>-T�� p?@��'����-�r>���e�r�;M�d�	Y�$D�8������U=,�A��[�p��	�n���c��y�w'�63��j��"E���{��������x�N�.��[P;��0�R�Nk�#?� g2X�?���	�d���y�(��ފ�'�#x��Sr̊�,�
��4V���$U���a�Z��>�u�ȱҾ�Z�ON�� �n�6
���Z�}��KF|k+Q|�@���e,n�^�v�����. ä���j�أDD�H  < �����,t`�X4B)���*���"���'m��l�^��V��|�kf�h�82V
m�ױ��ɻ?artŗ������s��L��R���=U_��
#�hbȃ��_V׮0r���9��[����=��n�;2�|��3D@�#
96`"⺡I#�X�0�0�Qȯ���B.������iȌ�7 �w�v�&϶p��9������d�����}@�����4O��(]*�J0��m��Zͭ��ɬ��%�