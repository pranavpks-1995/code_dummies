�aE��\����D����!�
gQ�5RM�a_i<s�M�3���G�ݯ���2
#7Pv��C��������!���ı)�&	�#4 D5��V�;�FE��L0��;&6��,�|U�lLd�0����X�m:vJ�F򚫎JX�s�}��(AUm��[ŏ|t;���R�c�������Oe�y}����Ξ��+���z�QL�@{��{:�K����٤?�Y��(  �!�ڒ�� �bV��XXq�U�"�c�a��{��?.$AJ��Jv瘃wa��ņ���_�io� '�`��uN��h�}���}	��l%9�s���fl�c��"�Yr���+��AjHZf'07@�� u���`j��+ªf��� &�0+�H�~��K{⫼t�c;�丷�   8!)��:��0��-d+DFc�����FU���x eJD"$��2Q�����Ō�{�ڗ�|�ě�3�P۾���_���o�ǈ~����@��f"���FAj����������m�,C�.%́d�L�E����4@[1hI<�xͿk���
`'�w���!  �phh�����zB����  !K�J3Z��:L�	/@mȁY��}��R\��"���y��9�0��d%�6J��ߒ3� �'M��W���Yx~�GҀs�Kk��)��eͼ)����B�H�8����p��t%,$���6�t� P�"��+`̋I��jpQx��#K8)��*Q� ��C�!��=�2����5�����1UN�E�4�H�  � �!y��5EQԄJ� � �1�\b��PY�Y�d"�����֣Z���5.w@2	��E�4�=�Q �����Չ� ����ϣ�:}y��Xh��6"fq�4��&������wuc��?f�82ōTT3�'ui���  L���r��CJ�I=�LV+K��w{���n>��0      C�u"��_� A� ��  @�*�YH��F��K�k��~f�oĔ�D��ˋk��W'e�j��+��%"�8Ș>�v����
��[B�h>�I
�9�Er$��U����%'�gr�m���4�'?�#����������_d�|~�gU`���D�o��W��� �z�@����8kO8�`%_�H6q� k#��Y���1�S�WSZ( w$A aY�'t«,��e<c	FD��� �a�!٠Kp)�*}7�e�fzO�w�_�_����D����+Kޓ�h���0����:�#(��[�D&�ݪ��X��DvAڔ�Ȃk�E����PƄ� ���º����~���P1�kdS��	� (��K��y)
��@�X�#���lZۂ�2����D���VW$o�s(�0�~�Q،�n}�W����V�f�7��r�g2'V)Ld �'E�U�r��5y�F�^�Z�q���s3E�����u�O#�e��(G��O�W��\hrt��.�f��i*~3�H��\��* �d����^�r�b�%���Y��H�Y��e��ӹNA�-Ö�0UD�]*�B�2p(S��-bs�����U�{ƚ�'�������#�3a���|���4�d�Y��9̦�����Wv��6�c�f��9���@��f�LBG���a�'L ��G���􉴙񳣃��aP�>&�Cn`^7$�JaS��]���V��0�`:,(_�Xyoh$��>I�Le-�<p�����uf���^J�8�Ϸh�Џ����2�mw�mW�2���T�Ϙ��L�D�b�w����oO����|��s�X���lc�G�l�y�&w�al���M��/�"P���&Q���<O��* �w�~tG�&0b��J���]�S����e�LPԶ
BɾG�o,���p��sR��{,Wa,U��O�U�܅A���v�ԙ�r��Mel$7�b �3�6Ul������	)c������k�L��n���í;7��`�I�ӳ�^�/���HfԪП������DpFz��]T(O���v��E�}>�/��^�(}��֢�!�k5]��Z�Qh�r��*�K���ʢ�
-9�b�߼�CQ��:�pD}��mrm/����EA��@�|�C�yR>����Y��/�A������9��uޮ@��;�����r�w��
5�����N��Z	����{ Ђg��dEE��eg�~tk�)ve��ji.���8Z��lU�냊��O��������D/{�jf	������b