�FU�[61'�ex�f\lªx#-��X���ウ��=�?����JyS����O��;IsE��򢵧�- j:e���>��v95`�3��T����+�9Y�-� -e��ˇà�%��1g�D5-��o����K�_�o�� L�� ����r�RD��dPNZ*��_%3��8��M��i���
 xg��9��I�K��axU�TV!Ivƣֿ���?C�%R,S<pWg2O��`| �á��� Because there are so many
terrible sights in this world.��
m�W	�`   �ȲUW�D:0Rb�q��캶�i~���F>��4 �o퓴�l�7y�?�QZ�u
��l�!L\қV�������\T��o��,Y����'H�����8�S����B��ͷ�m���p�_�����zz��\P�ĕ�����I�����qPlQXb��i�,CK DY��S\Y�	���'	zއ<��X��+�`�x}�)0��]x�ƅ�2F����z�\r�R�3M�}��J�B8A��Qw:*��+���Sv����p��\wC?�K;_m@*����c��1�цl�O�S�)���<bP-�جʗ��}�j/�-~�,���9���� �`���k�@�c|[��E,3c�7R2�8��dH%��iiec^�_�(EZ�X����4�����l���!���F������٪ �Xyh�Jr�J�B�3�����g��'��VE��۽kR��A��)w���1�����[�P��Ȃ��N��lwJ�̻#�M�\
�NF� %l��2�k�А��Q\���?��-�ਔ���~5g�26V�O1��	*^�*(�Ⲿ����7(���eu!3�ss�z�}������2�:���, ƨ�m$�Y��
^�52o`>�=��e�d�������I=�+oԊk�gPҚ{�	���/k%���c 2�w.IU�o���^�(r��3#H�H�D�s���V@5�@��*�<^�u�e�"�Ӧ���R�v��
���������r:���.����������/"���k�Wv���~Go�z��; y-x6<
�i�6Ow_����&u�iOU���e�|�9�p5��k�Cr8��������]���ߎ7��}�����S7��9� �ܷ��";��X����V5���1�H���z����Y��|Ҹ\�