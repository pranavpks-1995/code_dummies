���)��X)�6&��=bN��{��RQ�L�.���bnq^~��9up� "�#�e�����OΡ��I��"�pbQ��|�J�z�*��0�_���1��x��k�~Q�h��mv2M�+:)g�-���oa>����B�&���T��2�l�A��!   � �-W��Õ2=)�G��往�$~�L�e!A���X� !��PMކ��A��Xj`b���� T�5�2ڎ���5�г4�56:�Y�"D��Ѩ�2k�&.S��C�=Y�]�d@�E19����:O`�D�����n�N�U�y/�(%�O���<-�m� �s0�f���w�I���n����X���쾨��^7�(G4���N���`�]F���Yx6��t"��w��MV����iH� 1G|"nI>P�J��M�N�SO�XSLn��X���T�S���t?y_�+n,��^|�/��V߷?�Y��aL 9wy�u��2���Q�v����d�*W
�Y^/��_�%�
@fi|�R].b�8f�j�`�)�8ï����ڼ�H��x�h��r!%WO|:ϽH��%�h���V~/@�~�M�om�gj(am�G�e���:�s6�$i��Xc����ɏ#UWh��U���G$>xC�	뢲s�o|�EA�U���   ��h�UW�C��f0��oFr��öJ���3XZ�4ƫ�唌�Sfe��	�R*�],j������c�/wq�؅m����1Bٍ�]�P�F/�V>�w�!� ~�u|}�sUXtclR�
�O��T�SV��Uq�"Q	�(�#ŋ4C}0�-ƻ��%ƋKxe=,����
�=�vnC����2cO3iG�"H==�W�]!�M`/�&�c�X��P�����3�c��&5��AE�S���'�+!J7��s�7o������hm�������<��c�v��U���)z���K��V�J(���ԍCծ�.LY:Om�(�-@��?P���yԶ�A��Ҹ8n��:5�D��0t�� :�*�b��ƞ��H��Z2E�P��M3�h�3���F�T��Tg�R��]�b��o4�q�ϕ�G.�K5-$fl������M`Yj{Y���Ll�S*)d�*~*A�#ڬ�N=M����h��@dh�����G�ȕ3�B٩ݡW�(�p'7+�Dz���Ŏ!�{k�{|�Ҫf��㦠M�`ZIr�۲%�>%$<��L14����>���-y���%���>�H�������ӫ)uVr��̬8;��9<c���W�Bx��2@��9,�E�g�N�j �2�la��o�Ƶa���8Iy�B�k�JO 7��&�vG��X��b�OU��CN�&H3�!٫���͚9��l��4"A�ހ9���M�w9����x�$"�΍�
���L��0�i����6Ȣo��t�X	$k�ߢYk�l�LN�H ����g;v���<B�F�UY=�Uyom}�mQ��h�:)}����֟3j���<��7�l�;������v���q\F�������]1@}��%$
Q�����L�o��\��O�U_j�h���l	�;��Vq��{��E�B�m���ڣ?�y"��^8�];2˂�ʌ<�~I7�Y�ֺw�{��vKoF4*����p�{�6�! e0H�8e�:U�G�R��d�X�8f��5�Ӯ�M��[Kl��"lr�n{��~oq�c���h�o�6��q>c��Β>��60E��;�7�B����T=oIA�m|D���w�Bc��8��n��}z�M#��ߣ	ϳB�q���fH���r�\���خG]�P��O��M��NnL��OD/�p	i3���?D�f@���Abf+�>�X|'��x�ҹ�th޻ٛjl��\�q� N2���q��b*N=�]a4�-��ux��H)OH;��fD�v6�S�e��m�Cp��I�3��V?�������Qa���Kp�;�l�BT@}�J����U�Xb�S��4滕�����E2-�r�e-��*Y����l���^�����Q����+'K������dNU�����kH8դZ���l���<���W�2�#n��_T�}ͧk��]�^����b���-�.E㤳����ʦ_4�vp�K���abp(�&�_v;8��"n�B{�_?�Z`��|�M�M6�H�в�(C�����S1J�>���5Vt�:3��C���Ќ{���<��	����ޟI]�U��f+�VU���H�S5V�3�X�)�	���KƲX��cD�MV#��a`$(B?`�uP�R@4
~� ��}�'3��awe���Ѕ�kBp������\,�)��-�JL�C�^�����w����XFK���	Zb.��{ŃLh�ӈ�9����P�bN^�k�������h�������[�L�w�e/В�V�I���9�#Z�_C;��5�/%+q��D���\�lN�+�$�!����uo�����H�Yb�v22�ۺ
mŶ��X�D�������d�a��<��,0�2�}00�(���Z�ԣQ:�0=f�G��ǰ��^Rܤ��ǭ�:_)�w&�^�9o���m�E7u�.	�g&�ŝヒ	SJ�m�+�PN�ܸZ�Q�� �G���r�jX�!��[�1�J୾�2Y@G0��@L`�[M/��T#�,�?�f!�]Ю4I�:5_�nL�c[��g� �)��_�$Dw�x�%�� �`�A�2���<�!��������;-�P���ͧG�؝ZJӂo�*a._<7l�̮F���r��Z\�S
H}uԳJ�Y�t���$�=�-+� �	NM�L,�;�<