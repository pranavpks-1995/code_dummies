?[�e�ra]����q��ʵ�w�q���ci��+3��^d���\���L{)k�O�g *N
��)ݤ��\cE����Q�Ubn�@�x�����yI��䅻�I����js8�*���2�5H��ïˎ�R?�uw\�%��*ذ%�۳�ݪ*ib�ߐB����In�_��Wu%Qla�"ጯ\�my%@�K��SN1��p	_�B�u��>��.0��4c/��ߙ>b"�[�гJ7�æ�}�p+�ڞ�4���b������s�6-1F�i��Xar�j�N��^��H�G��iYR�$�L��P����j(E����K7Ip���J51�ej;2=��[�nm�˻��@﹢��F�8�pu��䪗���t�����T-8�*�Jeoea]��Kb�rҵ}L:�g�4�*���-����/Y*Y3(d~�S���n����q�_�Jt�To�j?��xk����!ߵM�@sz�hD<xH�=y15ƶ�r:b���e,e���;��v�&�i��K!"�r��x�[j^F�9F���%yA�:���x���B�3(��m�<2G��?p���NXKG䖷4w��r{�sw��˿sޙ���$�Q���=��5Qsja�<�^�ŶZ@����ԓ�����^M�o�~�./ɠ��'ñ'�����O[f��ʼ�3��e�=�G\�f�$��+�d���QY@d��Ev�i��k��e6r�^I!C�������9��?�bN�W8��8+�������X�~��tœ9f�0�I�AWo�G�2�8�_�����:�z��yAP2��s��ʤ5�k0��4�<�r�X�d�zx>\���a�ß";(V&���꡺�F��fz�Ѱ��!�h�M+=���Fky�63͖��dcX%�JA�-��Ae�t���6��ܟ�?���{�D�Ä�IXm�W�!����h�G�`2��B�V���a��*n�2�����v��}���Ri����v�;m/�u�@�K�,�Ő����-�6����(���#�\Ed�-���nw��dL!	�NuPo7˺!B[��إ�e8ח6Bo�|�@x5���˃�왑�w��~�ѥF������B�T�kB��lZ���񾃎��Vdw�lꪆ��z,Ug4U55'm����&O���'p��|�ƀ�`GMO���3��>� �(I��A�Go,�{�s+�"��@,˃�cF�fI��B9:�8��}�-��\6��2!��h].�p+��D�sn��N�[��ƒ!�E( Ȧ=��SC���y�I�<@1j��+L���r�1R�J��Pi����u�F�bBnE����f���\i����< ~��}�ߕ~���OB����4�u�gTI���7SA�~C,���#
���L �*.P�ID�����[UP�:s�mg�kխ�_n��#0g��l�h%�>�k��b`�d�=��þ�-4R�r����wK�<������n��G�Pٰ6�NB����f6#<9�R���%%=#��bL��%.W�BE5ŷ(�Y�q�ʹ[��5RgP��Tb�"r�_�����n��U��mՇ߁xA����!L�[t4(L�Ά�C�՟!iF��dN:�� �{���P�0�R]z���U ^�W"��k�m��+)z�}g=�4䈟����Ԥ�%�<_t�"K� U?%$������%c�V��� ��%#@%S���9ۚ��v��gi8oX\��+��]=�������um�mי��T��׽��Z����6�8}�V���79�,�o����=��4���5�2��G�Ս�Rh�?m��V�2ڮ��0�"��W���o��

�R�*����Ykk�W*O��M�d �n��7�K�5R(�<�9�!}�?����������rb�������۔Pt�Jъ&J�ʊ]��^�L�����JN�+%�[��~L6�`��� ]ȨC6Er��i��w)/�
�}q_k^�Cw&�3�B��0�g��!{���"7�gs�*��̒Z�Z�EO ��̌B#h\FХ��&�����@`����Jq2��m ��DXD��)�$ǋ���99��';��o�#uݵ���X�i5t��?174oVg-j���0G����8���m�6)B��m�x��.\�[�׾NEc�����A����
�x8�ci_�st2�Cw�'�p��F#�i�h�{�q&|��|L�?��+WB�����"�u�w�&�¥vOew]�J*������)��X-;>��b���	�W��fw��F�H=V�Bg��ō�YgD��,��!H�Ό4�ӗOVH?�(����7�0�;�2�!���{���@QQ-b���nPſ���a![.�_�t��w��p�io��u>cf�+�ET����@6NL��E���:�a�%�)�z�`I �͵�&;E��ɐw�]�tN�ŇAX���:m��?H 2R�!�����l�'�hyy��wDku,���t"�,ζ�&"�g��7�ort�MO2�RF�	�8
F`V���:?��/�g��P�u�t�K��QM��ؘc���8��;�����*Bf����c]������NP+[Ѻ�H`��/�zI��uŎuu