��&��KE��tӾ�$~�1L%	_W��o"t�z8w�N&4�M&*1Ʃ�K� ���3�\���X�N�ʍ��4X4�����X��);�琄�-�yǚ[��{_9l�TӀ �F[<؀�����#E " ���!UP���x2ֳ@!�� v?U9r �Б'�9ol���$���l�2�UD�����C"݌>
����*s�V
�� �0P��c�'ó��P���&�<��� �OV�p�����&i)D���9Rf1b�˂#��!URԲ�e�L !����N _圝�� 5�0Z���c5�.巭�p�2Z�s��!	�re!:i\K2B����$VDp�"��
Ŧ���I�� !ҁJ
���w���s�������y��a�3����ƈ��� 	��� �j�r�M�Bꥢk�A�� !����9�Q�s�}G�p[bũe�{m�a�����~:[�ݻtV)�<��A��@��T���{as�ł+Uh+,$8�$�������>_���]g<�`\0����N��N�~Ȣ5%4��}:Ol ^+�"����� �9*Rּ@`���K� �   ���K�c�D	☧l�*������Rg�iO!�8<��г�[�~��7�I���p�`����LBi���3v"mE���B�|B�P^��#]oK���"'���qֽU;��,U�a�����������r�����:�j�'�l�b�E�nb�!(yF���3�������]�ڒ��=�d(��̯�T�q�2ǭ�E�[���%FY@)��[jK��-�*�S����1CH�@�O���ଖ��d�=��0�WD֚}�q�M���H���p���ɢh����l���a�w����s>����E�h��V~���P]U���FG��Ý�iA�D�[,�&�/�/��O6�ΦO��N���ߝ�<W�7���f
LD?�����ښz�HV� 	� �U͘~��l����n��p\Q]J\�v�7kG2�������o���f���$)���&p������Pr�l��v��=E��m(�m�5�
m����|8 ��m������Bɯa�	�X�cd��E�r���Z
���d�Y�R48����<��bP6�}c:U�f�Y��,��ҍ� r��,ݲ��\�8N����NO�j��TɁ�>JQ��j?��c�7�$���oI�kX�P>*27M8NMg,Sb���G�zv���4j4���#$Ag��