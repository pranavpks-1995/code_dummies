6���s�~F;c9��.*��T��< \9Cw	1���Ž�2m�p�F�D�dc;nOÙn�C#��Ru�V��CW��Z�������\��r�E�lCk�6G@��w�:		K���R�-��B����6z|��QWþ��"©
���b#H��=�� ��w��oꉯ�F���S�	{� �5���H�U��p�"��܀y��D��1��h��)&kB$A7Y_ $���<�V4����y�N����6��L�* ׇ]�?��,?�����&�A���6����K�+���U��D�� �  x �F�U�$�N�,52#@ˌ��?�$��7�:�B^���.r�C��$��{��m�J!�[7�C�i�ُ%�����֫Kw3��瘩ug�<��_G�Ί��c��~�= 3d)w� ��#Ic�45>ɻD ^����$DL��%���Cqn8�<pe���{�.K�j�S�mg�������/��#�����ؗ�$W	A�ǋ��鴯t�Q�M�{ �_�g5~� ��k�~���o�Pm��+B�V���)��$�k���óm�s�B�(��?���SoC+�F�������4�Cy��]�?z�ηSF((��A�%7�(!�#�ԛ� ��d�}���ڑa�{6:uˇ�R뷥�k8R�bU��>*�ļ�xg�5�5h5���A�*�a�2�Q�jĂ�P sz�('��0�<�u^1�*p��~n5#A1P���
�|Uۻ���A���ԇ���8�K�,P��Nq���?���JN�
�Oz�	ˇ�X1��
��4��,R&�O������kv��d�F+�	9�Ɵ�AL�R�@w�#�g5�r`U�̄@�?G�Y'	�:��NDQ�B�ڥ� ����32�H8��֬8�
T�e�}K븯Zb�_����\�P2�וW�H��nm ���!*V ��ٚC��8,1h%e�ʔ�f�'D��s���D�V��M���RNEW1g�A�5��ɒNk6hdF4G�iS8a���\��4�'��Dt�{�0Ӎ�3�I���G���\2��
H�$�>�%r@p�?�9Y��^��)S!�-�RA��^�⹘��
�kP�'�܇�K��#��B|�Ĥ�\������	�E�z�I C�x�:���Q�B�����c<G��L��`W��
��K���jIՑ����"�5�q�7i��(�KӠ�ߤ_�/�P�=rpd�Lq�����P����ԙ��]b=f���BU��j�� �ˍ���i-��$ج�߆�<�_Ԕc(u�Ydi�٪�Ô�5tѕ\:�BZ�(�1y!B��R ����O��3}��.�(��U��|זq@~����Ō����]6�5�G�g����}�H'w#|�Ohp.���8�D�D��
o����w�O	i��Dm�$   e �f�u�  0���;S�h�VNy�C 5�Jp9
�^��(p5�-�jT������;�	����b�B�k3~��j���Q�x�@ G����I�-u9*�����J�Aw`(^30��:�d�ޛ��P�`� ��QrP8�@Z#R@���=�!X�Y��u��n`�N��}}�؈W��O�f�����@��n��G�y�A�mt8��
Ⱥ���0�͠T�۸�SeZݿ�j�;;�$�l�IrVR�\7 "Y?5*HA�+���~����>})�0Z��Jo���Q��3]�ƾ�,f�(pV�p�Wg�V9WO����M�l'0O�Hx��دr��<����x�6p^qI��B7��q���̽8c��fu\�;�'���89s�_�z,l�-�?ވ�T�\GT{iR���U�x��W�EN��]�ο�?�M=�#ݗY@�%�g9=eY1��Eu;ZN����"\W�Ў�eRb�/�.�Y�~�C}c�N~z%r{�*t�Z���e�bW���Z������-gr�@���x��Ȣ��p�t�rRߤ<a�#-�>7�������a
�r�+yx�
J���#�ݦ������)~LK'����P�������H�58''�g���w����Qb?LSMCJ����xdV�v^Ն�ʗ�^�@��vۣ@P�rB
P`<�oO4�'kװ5P{sW8���?�c&av(�|�DxB��̄A�&^�ǡbJ58�DtHV�K8,oN�b=X9�'(�Ѣ�#&�y��V�׳q���q�C�k���? sN/y]_�~g+8�4Qz+�F���s�MK��p�c9���0]���ޥs��nz�ԽZ8�NŊc+�6%+����I�5E�D�5�vٹ��.��%Zw ����:���F/l8�ܱ�|
N7���0%�͈�ÐK-�\�3�.ہڤG����r`���t-��3{ܗ�����v��0�Z� 
��^��"�l��7'�YZ����/�D�!3?)/H@`-+=eC	j�+����&b���+��:K�N�Cܕ̲���-3r@9����@	%u�4����T��Z-�jhп��(Z�yr��C��佴p��� ǎp���4sZ�(�_�@��CF�x   > �-������dL�V�%p½qG�YV� ���y�RI�r�;�-(m`������F?���*fa��|(B�T�t�aR�%�/��j�1m��O���jg*���~aH�>%�3=���P���=)*؃\�\��0�+RU(�/!-�t,�ꪆ�t�R��F,Я�ee�bO�qb��Eg��7w}I
��m������ь�rL�߽3J/<