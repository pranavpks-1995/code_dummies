����K�C�G�5~b7�K\��C�/O_�޻�v>���^���2�A����s��y0�I�zk�3Q�ty�C�E4gv��t�����r]��gߡE���Z��@��W�eFNZ��ӻ>���@Y�͂ [���5\�:l>��D�|A�g����Y����0P�U��^��xVA�D��E�,!%|�9: qWr���f���~|�˔��l� �r��ו���2�kT��g�#pgK�c�Ŷ���Xa�xѤJoGϷ��#.���
��oe�Iƚ+�»�<h��-�Fx�*(��֏�Λ��	��c�ƦXt
+�C��.|Q��nC@�X��ͮ�<2�{�x���^B6���f1W3ȹ��<5%�^��*z����}��s�S��?�(ڃ��;�y
o�_�~�0��*�: m���k��WZ���=`G�����¯������z�4s�G����<5�%���'�7���ْ����J���|5�����su���D�������/;�;��!��i�3`�%I�j�~�D��S�<*�4�ȝ�
�P�Jߥ��E	������;!��5��>O�w�§�Z��7K�����~c���v���X�ĳT($�U~ϲV��@���m�+΋@��({�}�#�jԊ̭�~��ۆ��BΝ�f����+��U���̮�X�`��z7�&���_� <U��6� pN�� ��J��MJ.�3Q
4�ؘ-7�Ӭ��Z�2z}I[�����!���5ȹ\�0ܸ"9�7X�M@�ΐ74�\���Q�'��!cI�ιR��c��0ߔ��)��F].���B��!�V憎��#Rt���-�}�U�m�C.3d���k�*���ŧ{����_x�q� �gy�h�}�����*�c3r����@i�
g4�yD�OP�Ⱥ�d��MAT�3� �t��]����e�{�˳�<���Ϝǣ����	X�uS��ȢQ�|�e ������n�tD��g���0�o��-a
��:韙$��-/��Yg\p��'H[(���(0}NY�d�۠�"���9�Z�5�@�AE����	{��F���eye�N�����E"W��q+���.N�T�,�43+[=LN�va2��q�초m��N�x!�~jE,;B���C���J�[.H��AkN��lQR���`㤺2�Sn��\�Yw�[�q^��e{
:��<���e����ܠ�7��䭎����A��-!Cg����f�`���G���c�U=����|�f�~{Mz��X
8�Q�E��1�EШ����ť��N>���Φ�#{Zczx�������*��R5��!��+����ғ��ԅ5Ȫ�!;V����M�Q��yv�[
`���mo�X>�0���r���թ��� �~��{�1Xv�)&_Tx����H�~�!7@�������g�Au��U���n�����e���C�lv�!Mm*�R a��u�^���W�f���s�
]�?�X�P+�U�$�5\]��˽������~�J��J�'����0�$����ֿΙ�|��s/%co��o~j�f" �_�#��Ho@O�i}>cb�0��)�#�No;�[���8�Xg�_-K[��8,��jM�|R��٫ԖyvD����O�[�4w�#N+3޸mgF��82���|'��� 뺮"����H`~:�6�_0���qv�Me�qt�V&�U��L8�߉��J��R����Vv�����4�-���Q�Q,�PG"\��{d�Cƌ�P_�!N0��>7�q��$OL�B���� 1���z�F~<'-�l�R*J��0H�Nf�z�=���!;SO3���Q�&P�/J|N)��ɀ#�N�K�Q�fv)T�T��Ogi�X���<w���<��e�-X
���'��@!�P>Y#/(FU.�
g�2��a��6.�xD%
d�`���3�h�\~(�O� ���lM�L ��8V#�a�i�H7XD/��v"�O�兢�n��-����4�ca:M��4�\�#+\?&b���T^b�� �)�{p�W��4r��C
��^;]���l�����@#V���E�<��.A���L?R�z���,i+�t��KUV��iA�'��e��pR�Dt�ҊF'F��Bi;�MU�g�����m�KD8�}�<�y��l�JWk�3 L�_��&c�N�^
�=q��-��	:^eϣIfIHP�=�g1����ad&�4�,�:�o���>����ϯv7oxo�O��뛳���0��T�$#E��?XI�N�j�*�xV8fͰñ��>�)&�-�����*���g�6�-e��b){V�1�a��S�cD ��M�[
��K_��Z�:"s�k��4��Uj�G��W�$[t�0�R���}�����|�x���D 5Й�h�>��w���T��3U�"�jTh8����;� ���i�4ꊥ��"���$&��p����~Z�����䅱w�
��{b�?��ƻ���'DiR�%�gě�=l��I96S5v!^��&���Z�XeV�f�^����c#����	�ڙw��?%�{q�62� k�Z27��i�I��3;-�I��N��a����(��k��cE��-k��v���k�)z�w�{����^�zF؅�[�O�U/�aA�l��t}��e��<+�j�t�9,3]�,�3>�'FM�q����-N���@��m��	Ȼ�Ţ���uR9Ux\��9?���D��!iս�
u���2�/�{U���b4Nm�x���D�fdLi|c�̳i�<�_w���cKj�@�!�L��c���sW���m��q�>�^RgSws��N���qwn)�b�I$a������,��D�4D9��2IZ�9��BrRy��nb��/3]&"6泍3���]W�������(���Y�Zy�J /��(�}�B����,{A�j��>F��jP����giO�?��E�}6��I
��n��{_Xig�n���+GU�.4׳�M�C�Ǩt��ʸ��������8�O1�[jJ��p��0c~8�q�C�
x� ��)��=2�\fh��Ӹ/΢К�=u�.O��a{�><��4�E�	�f�8��lN�}�%��`Rn]���!-��I5�Ye���VϨ�Bl����x������,�)}��'d#��j'�-[8ɜp������E"�����:=�= ٸ�GE1��N��l��|��A/RE���͔��JZh�,&���A��f�T�$ʛ�!j���}d��p�Y�_���4!P��CV�;���+�	�AQrwN�.@A��hɀ�λ��uWg5\z�`��0�bH}L�x�U5���ȉ���J�;u�vش����;訪��+��n�����A����a�HP����vh�y��E��V��k�g`Ui�Φ�m��0��(�!���~��E��N������yyލ�6���E��JP���2	��~.X�Kg�<|9�-��� �q4H5��!4C[�Z���� ;�ҍ�A�:�E8�W�c�Ϙ��$��{8�x��k�S��d2�韪�eE��9���S{Y��`=�Ů��A~t��j�!��g-���t���|j�������� Gh�4;�|1Biaa��^�&��^t�ތ�Kv/�p��#���?�[�/�0�![�KyE�g�R.H�����)�&R1��a��4-T��޽��T͊%ι.b]��_Vb�v��=8��6����w 
A��M^�u�������L��X@�[�A�_"�d�|�4A�Bd������d��le�{�6����� ��:< ������Z����������j��}rL�yD�� �2I��#"~��>E��ll��C�>�xu/��2�[��s��$!K�?��WL���pӆ�3i��"���ȼ��������K����*��$
�� 9t�@;q�}���!�5oQ���~�	F]�K;���c�
t'N�1r0�����~��-�w++����|�#�5��Y��#u�d��dЇ��^�H�*��.�5-�L*�^���aB�/�[�*_h}��K&���*EQ�4����=�N�w[��]*/��bZ��l���h�V�If΃��?����H�J/�l  
'��'RW�c�F�ؘ�\Q��P����P��B*�����g=��c��i ���v5_=��z���i��C3|7`��)$�W�ϩ�m�1�����m��Y#�J�����aBUA�9Z�����r��W2���֫��q���А��j�G�f� �����m�D ^�)i�8��0��?n�R�R�}��d��/�^�PDh��r��s>���ә,��nFr7X�‼��38�ʯˣ㯅�,�
���x�\�Z�%nr��᭿BvH���I*��?2\R_=��,�;����:PHvn8�6�	�K��R����Xa,�ku�>�̵5Ӽ���At��Cs�,a݌���L