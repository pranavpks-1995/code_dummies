package Acquisition;
	module program (Empty);
	endmodule
endpackage

