t^8[0FL�>W@�J�~d�0�!o�*昰�y�H��a;���*�����BS/���p���!U��\���Փ^CT���΋��{��t�-z����"��~%i'B>��/_�=��߄�l ;�V��m;n,��[���TEl�_\^	�o�I��:S�[P��L��;.<�Xj��	��MKW���	T��2f��z��]��:��1\8$p��M�&� r��Ǯ��������� ]_��p��PD�2 Wƍ�{��E6_5�+hN�1� ~D�*���������5J�#~���~F�w�O�fԾ+��x,�v��I�l�I�!�'�:ލ]]Y1�?[���L�l�A��i+0��������P�q>���jd�jٖ�����x����F<�O�U'J�&:(� =�$ݙ��<ۺ�:V�y/��Fa�$��Rn���F+i�4�k��VZ�n���h6�Y�Ϛ×�R;@���Ѳ�6Y�x��z�S��H@)�È}�Er>&��sv({'�%�j��-�OA�9����
px�\I��{���<��P�]�[�n���4ӵə4:.lgjm���h��K����OU����7���\]�n���0��w��L�IO��"����Fz�D��B���V��؟B��˅�Ѫ�vhV�I�;�tl�O~#oJ���i��43^��z�!?|�F�,l��v5�Ms� 	JW{�Elc��t$�jG�����i=TU����5 �F�97p�'St�ݣF�5�r�<n�s � \[�r���ɝ��W�`��d{�,o� �Ǚ���g/��Փ��Uï`��i͓4v�C�ϯ�Y?}^zW��|��Ck�ѯs�J8[��v�.����3�3<L��(����ʤ�k��^�f+n��&�H����W��\	4^��L��"�1���7��Faˉ_�h��6z��zV�m6K�
�.���s� x9֨�T���n}�U�d�Mc�(v�]������9F׫�f{�	C��ջ �>�y"0o�0
�EJ�p͹SN�{��nx���X��<p"X�aV��;r���c��ݢ���]D�C=ڪ��
E����U�'0蓚�0�2�s�ķ,/y�?h�9���v�����¯I<���˿<q�'xq�vQ�JtY�y"w����[v�fKs��>a� 2��B�/4���@EP>��
ih��K�z���+i�
�P�Y~N��&��C�T�%=ꣴ�?M��f��+�a
��ɬ�<���#t��Np	 ����kEg|��Qzݛp����ԃ��!B��?E����$�wEQ�ګW�x+N�X�
/0�s 2��[���U���ѳ5�1b<lY���F�����m��x��F�7����~��X��]�i�^m�;�My�_��\`�"���83��O3��Z}H�H�Q�� �_.��8�S���Zv�B�PI�S�A��a��ڠ�ʪq8�RT�zu-�l=B��/���L���R�U�}���Sp��+�7�FP0���@`�C�r��ɶ���l��d�1dY�!l��;&�&)鷀A���-r������
�ZQ�?c7H��Oi͘K�o1z��r�9}�,b���l��,�gߗ�