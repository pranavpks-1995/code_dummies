�F�Ѵj���Yn��b�*�j�����B����T*�g�	���C�|_��.���1ye|�F�f�!zN|��ܙ@  !��"�2 H6�V�I*�J���k��X�'�����O/��1Q|���q��hE3N�~ǀ�՘�0Z�/��ް
��eM�Ex�N����B��9�� �˞��'��FV�Ì��tL2�2��C�rј�6�P HQ֕n��.�	z)�jFTN�d�� L��`�C���Ǜv������L_��`@!���`�YtVg�� �+Z�v�^�(�S�6�O����/�KNZ�QJ<E��>
����<Hc%B�i��W��,��uZ�@A�J9�I���D�\���*G�y˻MaQ�R�_w�� ��L�U ���=�:F**W%^���4�����    !���
�a���N�u%K����[Z..�D]z��Q����iZ�U�:��y�;���E�5F��N�z�U��H��延$��� �;yr�������u�����驫����xD�Y�|�ps���
����>�ֈ�� �.��y˙s �!��Q�B�@�Yh��ËX-)��x���4 �Ȯ�f$O15���ύ2��<c!�(GSSk	#�.q\�o�U��F-
9�-:C��/ީ��>���lⲯ&v�>E'8�>C�w�y[Na����h�s�����