}	�.;O�����X�JH�v.K�TSnp].{j�mҕ^pPSLF�V0v���,�LX�'���$���M�"�<�,Gs_���.����s,LU�H��]XZ٬�\m���*�Q����G�濾B�������L]�Y~�� ��G�Q���#2��;7�Uo�m0-�2��5�#�t�q����>m��U�Qqv��S؏T�Ci@���2���\�Qh�C���VivْQ���I��C�&����h���O��B�7��t��NS����!�'�؍�9� S�1���sN�J|����ibR�X1&|�Z�%ț�	�8�{���Ⱦ!������@�	zek�xz�TcU?�D���gv4zX\��e,ăG���/����F<���lOI�tC�;�׊��e/a�S��^w�@h�BEy��U�$!�i����D	�c&��o���H�/�5��@W���0^!����J5N�߀��)�����lW_=�8�ibҀTo8.�6?!zd N�+�{*pZǴ�p�Dn�q.�������E6�̂�������!�{��;?vukc /��u�<� E�Χ�o�WP���"�Є
����1������hK�,��j����^PR� �-�@��j�
�x ��ûv�u�����G#���jغ�w�����QL�h�U� �" [��E�B1��9��t'$��*������J�6��EF�ag�� 8!�8��u[N�tr�=�X@���E�o���H&