	`6�9�.��9��� �^\	0�N������+l9�F��_d��,�� Y��WB��E )DD��~QƼԈ7��e�}k��5&@�y�hRG
^'ě���D�ήg���c�X��y���yH��$�k ��\��H�ȅj�i�`~.��E	n,fr1��u���\2x���b+�1�m�N��ϱN����$A�ȿ��e"<��J�Vfn�f��[������w����/�m�m�A.�æ_�&�2�9�}5�*@}�ܝ`(9g�Ϗ�A�դ�H�����5Uˀ��� Y%�b)�l��@�P�oh����v�fM���./0T.�M������oF&�!yk�=�,���>B�N�*�m�ȃg�	��u�U��4�xNKķb��9���*��_-�w�*��e�qn��p\�a�.QMX��:5<���m��
���Zb��]"�����:KVDD���7"��H�6)����WB���B������8�H�23�/�ˁhC�hG��+����Ν_K�,��!�F���>>�6P�=�3�����+T��[0Ӎ����Z��Hq���y$��=�)���7��ݢ���@�|��� !���6�<�̿!�aGP
��c����������쏒��1�9����\�@Vޤ�'S��^��h��;�� V���;��i '�qi&��m�	.�c*�S�	Ąz�ť��}����G: Z�~v�Nν{$��G��B[ �t#P]nb(P,>��'��@ 8�/|����j�"�N�i����� PĘÜ�7&3�&8�Td���POjqK�pc\7�ĪY�m;�$��B	�Z��^�>ރYX8;fB���o�]ꢉSNo��+b�0�Z-D�,ӣHt�g�䴙���B>��w�W�՞vR+{VR�a���#q2-��fhh{��X�k��C�YL�!n�MC�~zO&uB�d�JWG��I���K�J�HKn���|�N���|N4���Ll�5c,B�J��z���T�|)X��Y�,���޿����ʃtR��R1��b6Z��j��̳
�M�w��u�[�J}�G2�!�~�a�\F���ܡZ��"9��\<VFYXCc�Y���h|{p��Q���er��ڞ��mr�L.�Da�ڤt!�?�����-�9�u�=�C��\�M����Nh<�δ[x"��`p�9�L��J}@�j�߸)ΙS`LZ���_��3�2�#�L#�T�Ϋ��\�#w�ݠأ挰�kc����Ri�I���C�!_�