 	rv�k(fk�8y"�I5�����>t��a�K�����m~�͑�3�%쁸�(=��ӡ�uq��p�0T�"p�.)��s�d+�i����Z��X�����lF|;@�A�;$X?ܗ0^��tg_�4��*s�.��a�v�OO�X�JD���p�{�%r4Ư�b�ō��-�9F�Uq�r���uUQ��u�С,4p���D��bq����.>���;51V�������J2E��M5��{��v����g��.MCһT�����Ԝ���3ܱ����-yǪ|e~{�"�]���QPǯM�U�B�Ы.c6�C��F���*C�2K��{Hs���|X�>�쟽J<�:�Y&�_.f��R��R%Xy��D"3ۑ��ȫЯ��&�]���;d�.��Zۮle ��݈5*�?��x���>x��U�ߧ�i6w �q�f>��^bP~�@�������tYi(7���/�~5�ȏ��LZ����e�,��ݐn䬿�'����T�]��=]?�׭q�c�"-��x��:	�?8�)������:�_�YW��#ҹh�"Ĉ;�q���
�0�IƲAq�����Ц�o@Ybc�'��"x��^+�SxNp�?�i�į
"������O���!��o4`"��H�u�6��Îd�C\L>(�}��%��
��[}P4�I9y�x��/7� ���.��I�:�#<o����s�ۡѝ�R��,�<�n���uٕ����h�1۔�Ў������7��Kz.ٳ�6��j�YJ��Y ^�Ń�y�P��g.=���J)[�����L[͘i�jhtt;#$k���ۿ���,N�KI��p�&�Q�GFY ��)���_i�C�I_`��%:�5���(���x�j�x�i���,�q*�e�k�y��?�-9 �_�b���n�J8����V!ضS$D6E�!��0��ŕ���!V����Ä�	�a�r�í�"f��l~�Tgj��V|�<�Xǲ ����h���Mӱ;ĵ��+�0�-��o�� ��؋P��ƿRڊ3���?[��	��B�������]X�⊘�5���H˪�tf�#���r*�d�pq���x(��bz}��R�6��{ė׮�i-%�;ι�q�)�����T5x��8Tt������3�3�D7���%#v�H��{��_�4:�X���iޭ�F����T.�x������C2�/<	$K-��I��ܚ0"�P���bS��e1r�O��7��OzdO+��H.�Y�Lڏ�LLU�br/�Ӡ����r�Ö�ߒ����]2�Y�~�E���.�Y�V��x
�����v�z9�ED��c�K��J�R�zX��ǔҙ�ej|#�!��/�l����(|˗ ��h,��9�$����;� Q���V�s�y��7+��A�z^m���~_�����l����I��]èh��L�����"�,��R�͸�b�k�zZ>͛QH��M��|mm01�)v�T���z:��M�M���.P��<���<��~�F;�'�JA|��9n�!��!�*��|���\Ř��V���(��_ɔ�I��<�8(
��Z�����8mInaS�m]��R|F�e]'�;E@���"�q�����2����w��\k��* ��=�M1|#�^ ��qBb` ����-^Sp��T���^�؅-j%��