
(* synthesize *)  // generate code for mkFibOne
module mkFibOne();

  // TASK: implement Fibonacci circuit

  // HINT: use two registers to store fib(n) and fib(n-1)
  //       and one rule to compute fib(n+1)

endmodule: mkFibOne
