1�.@a�����@Q���a���o�[!bY�����!��;��#�w�3�7��Ze�c&t,YWR����Í~K>C��L� (n[�ج9�~R��e�! �%���{���.��d��o�P��8��~>����L�d��fCIO��`b�3ઋ>�+�zָCg�:t��q�0�����S�|�!hC��sd��C��@�:t���r��,��q8��4��i �3��
#`�7pfE��B�M6��SH��kš(��Z��U�ͱ2���>⫫��>'}@^���>�~�j�w;K��B�Vŵ�
Q)��G��Na@��9Ae�E�]�L��c�]�|;�Cρz   � �B-W����s
�JT$9�j��:�f 毺-g?�}�uap��C�PR�P��~_�]�Ɂ&���p��N%����e��(`Ow	�I0��S9 f�j��՘B��z��c�k~%8Q�F����N3�nO!�bo��O�[��˛��6�A1���Kn��b������Pǰ�^�G<ף�dd�D\�Kd�����n��{�,�ZTa�	�*ʙ���q4
*�a^Aȵ/x�y@��d�d�ũ�Ȳ�h�?��i�E�"���y:��Q�0��L������͛��2�o>@��x"�ٟ���ȷW6�W�4��CAs�!�1������Mn�3O�ܗ����z�e��<:���{Q�A�s	����4�O�C]����J��,���}~篖�Ė�� a��8��������@�
}\��uM��a��;�~0'�.��\�=A$umc,a!ŉ�ހVǋ�2%��Iw�`RY��d���Af��hɢ��87���^�m��6�A��IV��"1>���6c_�b`\���k��O��K��`���h���0G*h3�^]�vA�m�����Bub�y�7N'��3���r2�<f�|���Y�Z�?<��s��'��K�_*�X*����w�H↢��;��"��S�>��PI)��=>`�u�G�P}��C|�8�Kl�n����s�hb�^-~����RD��H��>�s�zv%�W:���փdf�{��}R��q��7F2<|���7∔�FZ���uu�ב��-�U^b�\��k��tf��_<�&M"4��Uk|�\Ό�A�Ҫ�����lG!�h�r>�]U�v�"y�FH�NV}�9��R{��<�b#��$=�߃ߡ������&�V���5x����f��������`�%L:P�l䂍3C8(��tl�����E{�}[����x�}߭���Ժ�I������TB��O?�!   7հ�U_q:0R|�0.��˙�az�p���T�T��{�w[��~d����I�ͺ��jJ����y���� 7�2�KT15��mn(g��0H����(b���$�I�+O�ʐCﳭ�g��%���v��-VU��Ō�4�����h|�z�2���/����*V��8v��7 ����@̪��x�cdk8��ѲVu�&�a� ��5Kޟ����l��P-���<?�!˚��'�DN��mg�NC`>rF�P���e���׀H���ח�c��W�>��a ��������?���9��/��BF�K�irz\�����f.��T�d�N|QF'�F��za���lF�'��`����	�y�
vd�u��hA��X����C�%�W�z�z<� ��\�	u�bk��^�}LF����^qG�Ы�QX���'ؠW-�\�6��