J!�V�����u����*��8PҰ��.b��P'�txE�ٗ�r��z�`Mz�)vAsޚ=.�6(@ 5����\�1��M �� @&m���ApA��Z�4A�^���V�:쎅�fS=�u�ͱ>���?���N�wK9�@� �E�s�$ ����0\�֝�b⒐�G1�a�Կ!��`�<h��M��zk	Ԓ;���:��⨲���B`f���6\��x���D�{NC��4pj��,<X55��<�Z��<�CĲE��8`�i�XM"Q�F��Ϲ	_c'ȥ������P9�¨[���o/�R^hT~3��G܄ a���j�������UuB"`��0�S����^�gE!n��]S�O��NO���'."��G����S^�ko�k��6,7�� )_xkkYb�jv�O���;�g��|�JR{t
�*EU�_�߯�P�yo��pZl@�֫{�'�󮃏%F�m���2ڠ�]si��$v�Z�K��V!�������z�sU�������/@j�IhEW:����X�;L[�| ����L������H  ��`�x��::��gF/�ϡ�d�ӎk:��}�]�1"��F���f6^d^�M{���/���u�.lLf�(j�i$c��jI�BG�z��D���&�!VG`���i��Й��ba:��K�!��mz�2 K�˼�LS�5��ۘ<J��J�b/z�'�%}�x�kv����?g�����?�I���y����}��[��qa������4�!2�?3s�@�Q˽_�w�3�p���B+��b��MA��)|���֨� �Q��"���h0��"�;�r�s�P�@��h����
'q<oM\ؿjD�P���2�H��Dj�0�u?��9�ϟ�£�s���v~�_�^׸����Q;&bc>V�c�w?P��$' �W�<үCXTH܊��ⵁ��˖hZ�?ƥx���u:򵜪kM�Н�E�|�}N�	�<��䞈i�+�<���;��G�*.G4�_�͈XH���d�p}��{���1V��ĝ-�%�̉4���ń>�f8�KҰ �@�ݱ<�@���e��f����&ph���
%�c`��=�F�
�5�"!��lc�"m�o���m,.�~�$�N�z���FrWLȖj�g=Rt:�&E�S�ʁLƶ�=I���K�њ�!hx|ҡ�EQ����y.i�o�rQ2���R*,u�xA!Ņu�^��&Z��\�ew���)$��x��s+v~"��NB� m�n�/b�/�r{.�#��+�͚�������9�m�8���E����ѷ�ps��$D�Y������8�7���p�-���Z	fz�k.�Ps����2ѥ1	�M�:��wc����BF�C����@�c�#*��3�+:Ȝ���{�2l#���az�d����;U噗�Og��$F�˫oQM&�Ҷ����$�����Ѧ%2
�c^ˈ��Eޕ0����ǔ1�j�ճ��2g<�5/�-���J`�Rѡ�/s{`j�o;[�#�,��i_���=�sL6=�m��Dd�3��n6�|���0}��t��Dd�B��خf���+��%��;�y�W9 UE�����T�5ώ��fqB<�L��)휠�tE�kx V���0�W��ڀ��b�7�1>C#��mhU�HoTK�_]��;)�^e�����L�Z �[����g�!���hp�ShP�Gb��FT����r�s�-E�=9b�<���&ć
���,�c��*��` �t�=a�hh�;��gC�o�4J7+�ؕ�,��K����w��{�må��J0�|��6駪��õ T����rCڢ�R��\�\�*�*km���Ȣ� 7��M�����ɼ}V��`r�����{&*�э�v�0���X���YJ��+�TG6H����5y� w�
@����Sn�ٹ�N'_`�b�׼�(�L��PIof�
H�R-� )yyj�[h�1H
-e��+�	`�#3��Wa��G߭|'C R��RʻaC[�R�����E�� ���Ҟ���!�����2�˼�!������[J9���Q?�4��b�St���0���i0���)+r�gP��*z����#��Ci���������g���%m�g�Ov��(��D��4(T�M{��E��ܥ�*��Л"��@Y���Ɓ=���v(C B� ��㨂C^����MY   !)��.
��APZ*s�*����9�����I`��-�r�����Z8[�gM'�H��m��j�0C��k���z�����<�Jd�����7�{~�]�X�*�axn%�A�J�P�
�O��Jur݋-5HJ�Q�<�:,��+,ΈҭA�<Z�J0��� U���1�HUR�ai���  !K�I4F1�EB��w+9%��Š��@h���֝�L-�:xP�{u��.����ͱ �r�����b�k|��S�?��<0�oA��J��lv|�O��e��>�6�����h`��X�ϟS�ɟ$�%��|�����-_�?�v�m�y[+ @ >�2����*��e/��>��M����4�J
���ĒDC��x
����|�3k�T��R�   �!y�.aU�TFQG2*��Z�G�#�-#9�{�Z,�j9�����R���~\ F������ #�[���4̺~��р j�;��F0q�]��0ǫ�����:����}�-N���9v�)T�p� |�xN��%j�h�u�O���~�D �   �!����E�²�
)� ��
T+:��&\���4q����Ƀ��P���ۀ�� wmFLk��;i�	���S5Ŭ&Q̧IʈJ,�NS��#!0_.q��eGN�*c���g9-]l�^����0����B@��7���~����W�_}�]T�    �!���T�p��L6�  �!Q��:��}��}������1WYt��]v o���{虰�U� ַ�  Po�g��K�j������1��ƪ���˴l[������U`�$hC�ݮ� CM�i�H|~���I��l��`B0Kv������o�^ 0 !����%!�h V �.�iK�+J��-�����I�9\��k�����w|�V<����Ѝ&�r:w�����ߵz!�c�K�q��KW�^�������lC�;{������-��Z��=#`��H�����A�+;f�}#U���wt���0�@    !)����!0��� �iWP�����"c�v�VcQK!I�-ڦ�lTt|0�*v)���"�u�~���v��F�q\ը\�[Bxb�OJ6<�ly<Z�E�X/�%�A�x1v��F�D��$>o���_]����_�)#����y���2D��7v�ۤ!����(�� ��S�� }   ��_�F:0Qd��M=�7os�^�����C��v�@e���[���}VuX&k;��"0Ü��.��
G��q������Q�kK
 �i�`���wY���6�Ia�m+����y-���E2^��΀�ǬIwU1 D.a� ߰��k��(��c�k_�@8'Fp����beQ�xc��� �"oӨ�wQ����軹9���*�H��a��<2����ޏ!�����)l%|���h^Afۄ���J�V m�Q\&��5R������N�m�s�??��m��j�9ӷ�2P�� ͛&{���mD҉�]�u](�΂Zm��4V�Q�]u�J�{�V�"�y����0RI�KA���"r�
�H���e� ��ٔ� ��E�k��CBA�ˈ��Z�iD�SnMb9�C�y~8���&���e gͽ�=���^��\\c��ba<n�Q�<R%����z����[�5	]�FpC�.���y ���45q�ebt4��EG��� M9#���sic+&}x�Hc��bu�*�spw�٤�v��E�_��=V)Ӎ2�7SG�}@���';h�u7�~at#)��u�����5.
�M�P��Z�r�����^�H�z�b�Xu`(bT� �&"{>k��ݗ�o�����=Cd�nq�������]�j �V���?N�B�!r�!�N�LpbD���,�5?@�ؐ(x�T8ۈ�j�����t��΍��?�$=�x��K�MÊ	S݂����f��,|Y%`�[���,��b'���\�ӕ ⬝�f�ַ��2{(&�S��\�ۻ#=�a.����B*��2��{,S)�� 8�ER񦯸q}0����q%�
�����M��l`���1��CŔ����>6�(��������?C�v!�={�����X*��*#���!)�4��D� ���e{�.�Xac���i�9��G�Q�1*�Z4r&A��u9m8?�Թ? S��ށ�<1߽�}�]�ե�c��Kߗ��-��&Ԙ���sb_�[��TE'O�w�T��b�t��U�A�>���W^����>U��C���	��\�;t��n��`�L֠��p����[1��ǯ4��Kq��'�ݲ�<Q�ٺ��3_*�PH- �_]D�~�-<���=��^s�m~Z�"����&�q�
�55�^w��i�6:U�Rp}���U����Ĝ�K�$z��a�>:�l������_^q�j���.P��3Y�M�߫������(�w�Ǳ&�}!/�YS�ƌD	���.�^���my��|�uт���c�S�t�&��Q6��b1n�ײ3$;�����E'e��2��&*��^�g��n;>�>���ު����)i6��6�4�����Ɗ0D"���@, �Z/X �A��Dswӥ�SQ}�����͎u����kqm�k}��\ʵ���񮽭m�V`mF��d<Y�y�5K}���j4+۞����SM��lH�N�[]�4O����{�8���K��-p��z�Hڞp����-{q1(��`7|Ry���峴�nʇ^2O����>|F籸Hx1ᦔ#K�X�އ��+��,q_j���;`��fff�2� ���`7����H���$p���wMOH������YM{VP�2��{�%�O�)�I�b��w�(*H�|����n�kTkj��.���a���Z��uK�A�}7*���$�)^�H�#?�S�1`�:�]2mp���x=i����<���Ƿ��\���8���*�=5���7;��,���B��>0)1#�/c�=E�KiQ�T��>�º!�����o�amhNʺ	��Z��(6sչ����N%9�濝��?}7ݦ��ߤ�z㪭��T m?��/7n��1�g�����I�nL�t���	.��3|�\�)O�<�;��&�d㋲�L�Nn��� �"\lD�k&�^���پCӘ��#{���G�.(tߗ�Ƣ\W������ut��fw���{���xˊK2.�ov�o&@EQ'I�~(xG������d��^�ͺ��!���Z��>��D��/���:2�K��	��ȣU�2�(��@��&·�*�X��?���`:8�J��X�;��M��b!w;�!�m�xUҶ6��{�)m�(;�핃�������/�f�կ#'�A���������߸`���̷���� s
=f�a`����
� �B"�;�b~2�K�+ffO��b8=��Y:.�'�Wv#
��L�Ƈ��ߺ�a�4*���>�W�d��]�Z(��C