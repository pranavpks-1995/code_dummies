JB��
��7��F���=�������z(��v)����$o5�h-?%}�E�K7rU��x��S���h��A��㊳T��6�$�e�Z��ѝ���Ӳ�M),Ý��0L�n��s�'+L��zUݱ�x��!������Āݻ��"�����E8�SH-��=��s��ZV2��ͬ��,
s��H�I@)4*#�2���]��`Sw��Sݔ�8�օ/m���}���,�l���_��&*�̂掏�_�v�9gj����${.�bz��`��-��:����������Ȃ# c� t|K'18��6}�&JN�]��^�K��fV�"�'��7�[!�^�X.����o����P@����]p�E8X�������~���^�Z۪��g�~M}x�-�Y�*����3#�̰�7���q�K)I>UL�!b���"�@��"`�x�tm4P���GX�\�@�@��q��{H �����؉��y��L/Xp���|�Mbn�;���p@'0�z��,�����H��:�bts�����N-.�h:9��Ԟ��l2Pw�f�s�8ys���w|/�K��≐��J�U���R���pc��sꨂ!0����}IU�):��O�
M+bo�&��eb��%���B��K��w>t��$��������'1-����2����IP�?A��y�JV��2-n