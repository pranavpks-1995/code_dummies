��X�ӂ:����7Zr��hCJ�C��M���v5�⛫����#�k��M0�O��aRy\N���X�ް�ݴ�]h��M}��m0���j�S�������5¯-E��麵Z<'I���|*]M�Ԏ�OO(��u}��,'Y^���t@^}����揯�����!�`��Oe62�Ƚ�6����&{L���g�	,)��m������%��D�V���+��ꚕ�#��a���tR���r,�2d��ӿ��ϜY� �|�?2���M���xx�?o��x=��b&C�0�:혬)5�@�˂{h�H���2�V�|��gp��5dPK:��O��u�0#���$�V-y�56�M��	S���wi�q�z0x�5�֭	3W���Y��ƽ�a�]�:b���ӾMM9'Ǌ��{p;��FΟK��Z~�0]8��w���ԫ���	H���V��L<�����J�[<��.��]5�'^�KG&.�C2�[f��I��.e�s�
҅3�qJ�g>8#�Ġ,���2Z/����EB�]��:�Y�u��u5�OHaD���k�7�G� e�v����)�
O�=ic�ֵt�Լ�Z�g0+���4�k��:ɱ�5�j#Ѣ(��՟��<��0���-tܮh:�&����mŏ�Qp�*v���"��,)��d��:���W~%L�ۈ��K�Zm�k�0�g�� �{D�[׭�����I��I��@K�����\LB�]���(7�7Q��
��A��������'o���8&��%
� ?��Lգ�)��D�(��*"���m��@2(���O��c��������w@�_��5��2�k��"����d�9�OO�|UƖ�i+��t]p��_h�Ho<{��+5��(�꡶>a<(�����^�$�U���xJ��߱T�B�(ٍC�c\�V�i���ݓ(�[\R��uh��!O�l&���8]�H��T�b�U����{���6� �<�at��Ú�������L<�yu�JE��I�� ��&���i|�!|X�Lǉ7�~��>.��B��N�h_�G|���w��t�o�1
���gU��Rz�!�G~��x�����i��8^(�RC�cA�4�<r�3��)=�3�Nc��w�_�^��-�h�@��Y�;�oU"���Q�ġD�̽d�Kl]���.2}9^�Q��
��SD�C���LV�����y)�q��[�G�_76��G1��*1*�f]��E51�5���$7�r}�;�����b_��(�v2d3��dE�Lt�].�\��`> ��Ch�j�Z���d��)�Q���.�&�g�LI��`�d���˟��|ԧ��.J�X׬uQ��c^�ln�0pc���"tMb���m<��Y��&��d�E1<Im~�h�"�fS<��kT�i���=���T������:ǫa��c6� ]��)m�G��Y)�ay�Q��o_p9���y���c�:"����� �L�ON?���u�j%~���?�5���0�[�}�Xa�尼�*��xR��*�|r]�F�����_Z���\a�>�� �OU
Mh5�o�˧Y�?� ��S������e� P*~�Dy��5�ͺEc�8U�"���^�j�/M_YK5!sގ ���y��;Hnpa���JL	�ј����.��@ʜl���	2�sY���aYY���z+v�P����z߂<6����D��/	@;��N��,qNd��F��P���.�ܡ�˳r��B���#O�ξP��lȖ�n��|��F�Exsңrx��`��:b%��as��5
���p����Ui_+�����3ÐU�_gf������9�B{�ަ���ŭK�f
9��b�U\�xF:T��v�S���O"f���AY�w���uǻ�~��U�\�tZF7��"�˙��6��Q2�~O����%	|	�u[3�=�y{�@֦�;�$��¯ocZ[�F�{T
��'�.)ǂ5ב
���GJ|�(�j�T#�?F_b{�������5�>��|I3��n|�?�-=�z�4>@��"O��RY��O�/X~�:��#��"wl��6�q}r�$ѳ��o7<XI� l}�{/2�Z%a�G����t"�.���~0���*�Y��-�!����Kt���OC��B�~AX�P\N��z��J�"�`8U/Ir9��,PY�`�v��_�MP��X������e�cq��*��C�_|:Du(聛a�wE��]�|��h4Ż^ڈI��'�_k�Tċ��fw�(6�;����pZ-DV��T���pZ|�zKU���_�l�a<�4Vh4u��M���n�
��pWm�O)E�d��Cf���<��7���C�R�~Y.5i�������/���n"�e��&x�]���7�`�V� �C��Ci���W��/��?��3��7�e�{�v����0T��@��Ŗ��mÊ~ء+���P}���~�ns�jAQAĕA�P�K�m��}�%�*�$lw C����-�%��Sږl���/�.�o�7Ϣ�jƁ`N��/W&g��]{��ݥa����\�#�6����z��]w��V���])k�F�Sf��ތ����$���~(��=f�&J�4F�r�<Π�~7����O1�����nd{��N�'���Nbzr�Qk-۷�HߑQ�AZ�����ə�x|�%4�3O�U}��MO�p�kf�e��\�]��園ex@�,Zz#�ʅ��Z��[/[���۳Kx�Fn~K��kur�k�/g��pVmSW�7%�۽���;�$�ľ�܉�Ϥ
�������`��Aq�d�t���tn0B0
R����&�I�cAi�J��t��%��ZpX���T�C��(�[���$Tj���,�R�n��F��N�)���h��%�>
E�J��oJ�Z�Lҩ9X����-��9qص}nN��FNx"��N`T x%|N��%EVƎ���qq" U�j�]���G�s�$4!��h�4q����-�P`ĺ%9bB���_�����<zJ����#�:���!��3~�����K�p��f�O�m���C���(u�1?w~nx�0���s�1P�r��/2�p��Ș*����6�D&�T�	��P�HM3�_H�C�>���i|[*:k����%=�B=��˴TGg�y0�Ujh�H;����/�<a�R�"��UZ�[���< �`א�>E|K�y����tSM~�״�0�����IcfX�ʹ���&eУ˶ӛ�1��R�KgE�IF�/�3I���^e���G��[�M��:�\���^�DR�.�N�t���-=���ߨB��o�[c�]��	�\�)��w$�H��a�����+�s���b=���݃��$I0�2�����j�PS�T�~���O �_"Oy* �: f}�������"B> ��mXml7�]���
8.��I�K�Y�\��P2��_K}A�2�n�1��s:l�̵�@X�2 ��UVy�s�� ~����ݖK,d����S���%bݓ�3Qy���E���̇?`&��z���;��`��������@���Ț��(�ХW2��q ��n�d�0�	iI �j�?�њ�o��LWH���;ڕ0(�=4lǓ�n+� ��;Ȑ�s�NS,�~�� ��t���E���L��:Ʋ�H�N�w{��B���^��w�I��
u���v|�6��;cn��AI㧨%�3����엩���Iv����%h7���{�n��-kE $NNN��;�d(ӑ���B|���)��:�-��W�A� ����Ib�BVA/�!��Qy���_:�l�����Z��5�o~e��h8vA�믦�E�����^H���O��**+ڛ��N�K�W�N��RW#{�5i�맊�1�I��M��e�j�!~��*�D��Viy���:DTOh#�����_g8��6�=tCL|�	�D��'��J�#o:��Q-��������%�D8%�³�~�|M���G�"�a�W�
����jkS�}�As��K��!Q�?W��~��b͍3z�
%P��V���.L	:
�����7Jϕ���Q�v����F��B�5L��Z��z���C�s�����F�Pa��w9�V����iA�E�nq)�D�7�$l��_�|�9�=Ű�4�m���|އ��	����/mKE� *���S,Z��ݒR-!�c�^i�B	�����}���H�g"��C�&�&�v *�D1}=QB���Y���ʵE��Қ*�+y�/��D���sb@�>��:hi��Ŋ>$���}��*����n7��ZUt�,���$���.Qfu��z�@Sf��?HOk9�/q�VwS�3���yG��$�Ho(����