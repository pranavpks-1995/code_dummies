package Lock_Detectors;
	module program (Empty);
	endmodule
endpackage