package Acquisition;
	import Initial_Settings :: *;
	import Real :: *;

	function Result1 mkAcquisition(UInt#(32) PN_no, UInt#(32) ref_code_raw,trackResults,settings,rawdata,loopcnt,channelNr,status );

	endfunction : function

endpackage: Acquisition