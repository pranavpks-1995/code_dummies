�ZP[���za�x�t��o)����Z���F:���ⱍl4	׃�Z������J`�&�#xfH��8�8��x��
0��*8R�pg�� �B����*�Aɧ&�b�ZP�	b!�$F�t��>=FA�]��!�ӄB�MXރ�=�a:ܞ�G�B��scbj��F����~�{SV8r�L��O��9�<u�"�����&�A��Έy�@�S���}�,Z.��V���9;�J��w}	V��v���H�J$�y ډ�"���03��V��T��1:�@Qe��兲`A7�Z)�v:�������,�2K,�����&Y�#����V5���C��l$���/��);R(E��!�2Akz��尿����:�0��PȔe@r3�����5���	��e �b���w��I�Q�T�oz�l$EPz���b��X~T���7�׹���u�daH9���Jj��v��r������
�;�乌�$$jv��	��i� 7�5�R!��V{@�w�Bc�t�c����MX�����Ƙ(a*��C0ӎ�9���Y�Ҩ�u,��7��0Q�g ��D����͓��p�C4�ē�C9���و�*lx��g���N$�������|����y;�8��-�Fq�(z��:�Ȁ"��L&��ɾ�u9~ʌ3�k�����9Ys`�<=3����"��8g>^�R�/�
�>���YJ�|�F�{���cZ�1���M�ހ�D2��   * �B-����!"c�/7��Џ�$:�f�����,��rA�h�/�V���"
�0�tY�*��Q��;�!���
iy��$5�fP��W�%	)k�`i��Y�٦��I�F��7�t���A0K9)T�@��IIU#�?���R�'�\2���R/�sC4P���S�fb�ӂ��f��{0
kT��Ck{"���*F�ZW�и����L[��#7Mw+�� 7Ijޓq�T�5���MACyr�I^��d���!s񯡚�,�F�mj*O�hN?�C��/����p�f�H�u�e�1������6�5Wz8��s�5�R,K��&�e_k6���ÅHQN�H/=�e**g�A��a���`
�5vh�մ�S�	�
��SB1�ic�4} �����P�k���������j<���ꝙ�L:�[�6g��[���T�:k.�/�)tt-1	����>
H�$_W�ߢ����G=��W?����&-I"�g����s��ei��3�'��������%0�n�	:��؀D�8Ԭc�g��9.-K5�ބ��-�G�ךH�
p8��.׎Q��B�6����1�yV�I�lG1�((6�|���fE�ȕ��!�|!	��5��㈼v�L�YZ7�t=�A)R�
S�!�p��cRj�3~ӱ}
�ۖ��i�vfY����{.d_�d�&~�!���J�䡣G�������G���IIcjv�@ �8������ص_�አ�z��ո�n�ƦO��Lݞ��	o���U��a�b�:(��! (�0*��#�O�w��{�*��V�6����
��?6�vַԁZ'�8��'��v�ŕw�ڎ&DO�`�8�g�*V��0`H���rҶ-�8�(=����OͶfJ��Ӕ�j�=Jwom�&�4Y�Y?�Pw�ц�x.�Q�uD,�`�F���_����ryWų��Gl��#�*89I�y�ne�g�����sЄk���^�|)v?DBf�� ��ʦH?�G\� �,��)+�~X�B#�^���_�p٣S\�`XD���Q�0���ס$U�,�/h�El�	z��������!����ƃ!`l��(�@��gM��A�#�>��yI� <��sKv�,a0P��2sv��O2t��eʛ��Tcv��ɉ:-P���)	�!��[�Q�dO�2U)K{�ɇ�V�A�#��TC��Zx��d�C/�P�S�E��嶁$̺̏N5i�Ӝ�H� �����US�E鵽��t�    8!����6(Pl!��  �6x�8l��F�fdb��N3#���n�P������Ʌe�P�sF��h�T��biu��o�F�h�����������ڡ�U+B�{�I.ѭb���5k��� <�pu��t��S;y����޽�np     8!���#�	\l1F�Aaǋ 4-	�:�^��1��)��)�Na>���|,���%��.�����gs�G��lj2���ۆ��o߁���%y�xL�^��w}���(~8L$j�.��LفG#�� +�`����Ξ�P�%�A� y�H���B
��o+[�@`  !����30�b �����d�������@�B��~g��j����	�����U��rժ���/}���kU�k������c���Mh�����ΚC����U/R�n-�k)Ҙ ���r� �@��-/�$�U?ݷ��oԏ����=;��� `    �!����� " ��n�,|il)��8�u�=��P���]��`��S��;�}#�=僫�8P�F-�R�Hc	4�/������8��4���>m�w
�k�Ki�[�o8�[��
�2�	q|�l)��8��x^�cwT��/����w}�����    !���b��hP�9��V[�·��"�(E�����}�9 �CӿL����K�`�\�������̈U���j�K(�\س�W�F�ޞ���Av�[�V+�In�>(�`��� �"�J[R>�ݼgw�I��UT�����������1�ݮ�n���yۛwP !���C�$