��C� z�T�-sK�ٟ�C�1����?%d͸�քX6]uB��m��ۚ��3�g�!;�>_G�E�Mw0�a�1ϷlѶ�r`(���f���o��uݲ� F�bY�J��o�)�3[U�u�K@�|�
:�y)\��9qy�S:�>	������Z�����!�����k@����������p
v�݄�5ڞl��\�S�po�	�%b�	^�Fx��=�'g�á3!U׎7����MJM�qQ�@Xi.�2f�����
�+�X�VW[6�%�$�T;�:����A��;"�N�>
h�����G�&R���l3�BaC�[A�Yɦ�ޞ;ѷ����U�)ؚ0*cDD紕JC1^#�|I������tx3T�g��Cy���v���_���q>�q��z=xr�'����/ �Ge �y�7�x���g"�^P�ܘ�P�*!� �����:��r��M�c��c����oW���6!ȝ�)�T����qe�m+��I&ц�	br�h�X�]?14�6�!��8y�H�-�Sȏ��X/$�U����ܖ�N3�K�eOHn�n��r��1�sr-���� 8�h�)�[�E�c��!M�þ!Qz��7_�A���jħ��w�e�1f���lz���e`KͲ@_���&���.91k�oP�Ȑ�s��DG�lB��2�JXc����R�R_g����]#����K<�p��q�TRC�������ѕ ��7��"+1Te�LQ�<j�a��v��a�@�9���&�0���Gi�v�#�0���ʰH1�����J!�
����-+`w��d=s\�b:K��y��[ �?۝��t��r�'T���V��q׈U,W�����˹����q��Dѽ�޿�G���93O�l��F�\|_��X�rqG��k��@Yo����Lu(�p��ݺ��[��Ե��ˌ�ߚ˛iP��8��g��PǑ��\j݆Mx7=>7C=�N�͕��y�r�U�TƂ5�_�!:8��j�_�8j+Ci�V�ïs3����e�p���!V�k�5�8Wg�)� �����Ƽ�M��Y�&�5��Ǒ��G70�E[r)z�@(}���9r7U�w��
L�#���/6v��(KM�7s=���B ҩ�!J	&/.�3�4���ʺ; �Y� � �{�Wg2H��I���,0 ���&][�Q̾���|�_�;/	�5F�<*�.�����,DP��/��ey�5�..T���| 