�M�>A��W�E�M�%����� +DtR��/K�GW��Wڄ<9��P���,E�~d�eE�9r�����v�C=�ӯiŮ�����*O^@B��fJ�+�	S��.ĳ:� {H=����' G��^�_�א�!O�)�(~��jwL�����0K'��% &0:�k.��	^��֮�^����z�L$pe��ħ��r~�x�ͣ�)!�ś��k:��Z�>G,2Er"Iq�J�mkB�D,�MV�H�jM\2I����H��,!�;d5���� �6 G���U3yK@tS���kTJC���� <�o?$�h�5A�)��,�Ӧ�I��v�3򤉓ּ@.~Lη�,�}�k�|?��9: 9�A�W1go59L�/�{2��[�k��/W�aM���7'�W�?�y�g?p�i�ʎ�������`b����Zg�_��YxNRA�'��++o���z�#�/���=��׃C�(�̈�u��a��Ε������:�C�	ۨ����{�u�� Qn�)���3�y.2,��?��_�p� {���p�n܅�\P��pC��w�'L2�F>7��>���A��G.@ e]��]똆r�o�_	�_���@ �l@�K�*H,_qM��o�X� ;�$]���h��fXF��b괇�Dj龰�{/�����L�F�6�
�������J�{r��jD�(�I���A�����r@����+���^�
�+��gI���顢=��[�(�գ�J�}������J��E�v' Pd���\;��<��t�2�Ȋk_�M^歶��Ҕ��]Z�����mĵ�*2v,����C��TBf�T�|G��V�1��s��N"蔧W�{s(��6�+,������_�v����5��P��Ke���N��rYX�/�g���t�eɆ�;�q�ܳuȊ�����p��3�?����H��[��F�w#�1�Ǭ�~���߃�V��dm�kd��,������޽��(�a�~hS^�P�oPw�����O�^�Z��_"�*zx��
\?3$�А�&��"샘N$��rO⵰�܎��~0�]���ܓA�#�h���岞�?_uP�=���&`��?_�g�k��4�VY�a��V�2Ƈ牻抄M~�a���GƱQmy���5/xō(�C��Hr��
od$Ρ���Z���y����
�2����x=��6�v�K(��zcTP�B�;wǇ�rh����,f�};��zs�w�V:両�!D�5+��p�*�'����>��\����3�01�����d���٣	���lD2�gIxi���\6��y�6��� )
���z+_O��~kѐU��*��Uk��wfj���/��c)Ы�r�;��GK�u��bXL8 �u�Dy?�N��*�����%�1S$"	F>`�p�:�<-g�!�`�������M�Orг���C����T��I�b�:���ڛ���φp<�]Z��*����U:��2��d~��l��o,��)ӌd�3J����I��*�Cg��]E?7������E��R{�Oo�w��}\�|A���|��da���u���狨f��0ޕ7�n��v�ސ�N��ف�1B�Xe�d���--��y
��4�e�����y�@����b5-	����c�^4�=�y�=L��O/��o�p�݁��u?-ܛ��3�>k���������[9����7�gK�Ǻc
q`�:>|?/^����*�+Kn�"Z��;)��D\[^