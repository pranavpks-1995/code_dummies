�^ͺ�o��h�+�R�TJԨ7]3{Ꙋ��}��W�P��]��f,D��y��w���pAs�v<�(J쥼�h�W;S��KX�v̌,��t�i�'�� ��#���h(q�*��h�����u��ܻ�M춎1;�3��TF���;@�D��   	�x�W_q����H�&ƆEd���V�MnLkʗ�������	�4P���[����Ɲ�Ww����n��+� pZ�)�<��]]Y[|�}"�A�yD��͆�:Rg�O�)�)�'I�XW0SpZ�a:j��8��*Km�	�J2��̈́JHs�Uf���G7Kˢ>�5̒���)�7^#�5�/��>��_qhp�����ְ�_��:�!ib���=R@�W,�I*(��A��*6M���1��E��٤O��K���yN�����sp��ۑq�Y���]�&�ߓ���͞V8�O�S�R
�Tq�Rk_�ˑ8��d;%�����ο�sm��d�I-a4f�+��� ������������s��Z���Y�^=�]��.y:�% pv�V��/�w��:�:�T�R����ORĜ��|9�4�;�Ut	����>��B�rh����D����LĔ �x���^.����I]�$춪�.��1.K5���s�������`�k,j��;"��)�Gu�ִa�y�F6�#ߺ�����!�j����s���r�P�mp)�,��_��4{�$�d���{��a�g[O���F���y}9�3�å��Ho��+�V���P�PZ&��6FW��r��j�dW����h��i�zH�8;d�4��Zl�>�m3��"2�����峐����+с"�&��*�}�b��	� e��a-k�}33m�7��j���lm�%�-�p��
��2�@12ԖM��Gք��}��!����\�B�7*.�I�H��!�	�ţ�a���6$F`��l[b3��?G��m6������([D����C��x@�����!ڡ������)���[��Q�c�I��[cۤ�<3���P�nkQBNgV]Lf́1:4{�8��s	��c�5s��Z�T$���9��WF��n��*:����hP�]_1� ���y8Hg��:@��}<5�ێ<��E��{�J�ؗ,Q�c�|d�M�S�\��`�AR��  J ��-K��:0��T��$B���㠪z9��~l�ߓzM'PG�;+~K.@�@A��#��l+��|:�NPӷ����'ST[�O��f�l�t���<�u+Ӣ�9}��$���_J�H�B�57��5t��W�l�Y�_n��q��v�>�	O�Q�Q5�fp^C���� ^K���N�";�K)e�q�P0(�U���hpD�C�t帓����ʑ|��B��E{����c�������y.���b�bBe��(\�jSh�]�Q�@�v	��NN�*bխF;fW�?�t�%��̝�E��N�������K�_uS�@��]� n�p9�C�u!µ��� S�  �  S*