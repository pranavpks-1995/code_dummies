�$�kX8�'pRȠ窰�N��-����G&""�T<��� o^�b���������;����Y� �
׊P�I7YJ�S:ِo���e�m?�0�{���p�<�u����C�9�����:KS}r4���C��DD�Ei��������-�>�О��=w���}�{@�P��r��[*-�'1�����h���L����?�a��7>�p%P��L.-�$��=���n�V�ؖ�6���9�z o�}�F��9���B1x~
���Zx!��4P��&��z�>��q�Ů~y�Qsb
o�����14�~Oa%�sΉ��r�6�_��m�Q9p���}C� ޭ�3GvNCa����ZǠݽOQ�q���}
ۄ����I*��F~���h-ٰ���j3����a�o�k�?_H2d���y��
-SPi�1�m��_��3�)�z4\��M"��� ��[;?ў��95�~��W?.�1y�dv�K4�7���K�\�����$=�p�M�{�cxrrP��Y�0w����}wqX��80���2��H�Mrê%Hg�WaЄ0��C9��   1 ���u�|���CnD6,�@�T�,^h��K�
g���ʌ"L�����O�p�S2$^�i�����������'��U��^� g��{�lHp��g����x���I�t1N�ͣKX�`�B\OA�/���=��� ݿ�c̢l� $jh@���c�*yS'��o8��v#@��LSn>dd��`����0n���ø:jC&��gj��We���ДU��98�li��;���I�V"8�����UR0���l�q��\�w�juӾ��1Ԗ�'�4���p @T�P����LR����wG#�eJ2*$Ζ���6�'�qt�6�ҁ����ti�����&	�O�pI��Do�#*XT��⿌@����A�:8p^@z��/��KD�h�R]��m��d
�1(8����a��?A�Z�t=:R����utzd�]mE����3���v��@��Xɧ�+���Wb��%]�������l?��M�뫾����;���a����Nn0p1�MaQ�t��YL�ɤcO>�2�ŦEr;37�w�}��MGKb�\��_E�ɜ�egv����]ˮh�6�C��] ?B����,�ny�+��V8�6�PcI�aode��:@S^r�Wt���iX�+�����6��<V�Ls�M8'�{'�N� �}����V�z�b1����-��.٫����5��H��ד)���-�A'@
/ ���J��~�I"k�\��q��ȁ~FM@	h��YD��/��x�AV+#Cf[� _{��3���ϟ����(�L3��/���I�]�~����Y/f�1)iD�(��(��<��H�B7��   / �-���ÿ`��uo2V���&��n�;��QОhB�r4���.���k]��� ��fL�ۯ�oo�� �S�e	!_�t�x�"<E9� �|Rc�p<�Z~,�����twڴ�/@шVK�>	���?�",G�Ú�T_ķ�\��ʀ�!F|��X���y�� 3�H&�l�Ľ���A/4�zL�Q�}T�:t�!.(:k��Y��5�Jm7'U�1B:(�娈��I�W���u�pi^3�Uv���U��B��|����ԡa�F0Jb�3J�œO��������,Rj�c����}��ٍyo�ǧ��T��e���U��HH5�x�Z�٫9���@�6SCG�ټ���&j��_���䧧	�z���P�ECBu�4�n����auI���P�]�E� ���ڤ�2�SО��8�^ۋό��"	e�D��	S����ф�A��I��teU��I�e9��^�mY�,>�8�2�`�-������Fy���ℜ��j�d�,8X��T:��q�E�A�+�)�~X��vF����̪Y���N���   ��p����D:0M�Al�;�z�ձ�����s%�~w�6 ,p���)��u��*\��<������1e��j�4mY&d�F76�����J`��u�5�F[.�h�L�K�ÁG$p��/���/� �
&�'"���C���b�8�X�sc�U:�+O�3iu�Q�[窀�6qK$'q�߃ �B�y`aX0sgX�����7�<X?t&�=�`�������ܱ��O���D��t�>������c�hJ�MV~?͊5r�{KP7c�Ń�ћ�s��U r�o�eR3�G*h�� x�?�vV�"����z�
�._�+!A�w���P?]�r�|g�>&R26�������i7RЩ�`���,�Z)��:���.���