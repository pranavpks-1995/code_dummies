�~��u��m���p]+�ϖ���h���B������2^|�$/���r�\�x*�ۼ�Ohc�X_���O�RA܌Q���;&��<�W�i
�~1`�bg.��@�}ެ� J}>��^��?��*�FJ����-�M�z�P�ծ\&��Uxx�>���y|�� C��$�S*�=�n~�
=[� �l�ӛy��\j���=<�������T��˺\ n���@)���V�������=qRd@�u�1����@�҅�+㼳�r�l���WU,D2]�����ɠ�g�t&����z�Y��E =EHc�bd�\��,�苳'�=����PIr�IA@���n��o�J��]�V.�z�)�'�Q���V\.6�2�5
�7j���˙�-$�ʳhX����u]�<i�\u�S��d��t*��\�k��<��vk�{� �˭r=�\b�
[����CjT�ׯ�]���-�o���|��;Q���m��Y5�_�V�	�?�5?�Pܯ���
?���k9�x�JK�Xڿ��\f�=2�H��	�����tG��_�6W�+gYx=���s�yכ.����di��"�h�;���V.pثO+x���㡴U���j�=���R�O쉹~�e�A\�1�KdQ9���񀤲d��`��H8�H!�X;�fP4�ƣ�e=R8�O�NN�4}�&�8xF�
``<��9tu�T��O�X3�i*���QzftT�+��"N��	|p�]�ХQf2��hհd�%�]-��Nt�؆L�0ޠ9��L~���h��U_`�|{�z�<˚)�|�
#�!e__���g`��2��2%y�7���������T���d.{8��r����Jvx�§�	)�
���G�n^)C�zW��Y ۧ 0���u7�����/��+03m�MD�Τ�+	cMR*�O��#�$�0!���dDYG����~��~�ϫ"H��c��E� �s\J9@u�e�Bqm�&�mI'�#�?iQ�)�X������:z��0�@D6dۼТmx���A��ؑ���8�!1e�,-Y�N��0�?�CC`Њ3�"�8��CTl�P�����R����ٔ�^���3���Ʃkh8m_�c�-BQ�<\���]Q�$e8%\AUƪq�`G̐���v ���˅��3!��;��ӻ�G�/���GF�.�?�T8�qE|
�{n\c3R���3}ϔ���
��N�J�p����;�A�B�!����C}W����g�����Fu)QM�B^«�D�1|��g;��dci�d���Tv�dF�W������0�2,�؄�>!��m+�Vg�'�P�?��pHy�� YIʼ(�*��Vtz�WThՑSV�K6�-:N'���ϗ3�
�U���'�}bɚ���>
�����6����O\iK�-��){A�$�Ɔ�t)�r����pI�b,1�Ғ"'�1a�B4���ԅtD��1B6'��qo��I�R�`��+�)˱:QQv�$/����z?�77����38�=IM�aƙ1��c����o�s�}/�砍a"�\KF��
���v���� �~T�57�?hݙ��݈�� ���n�GȊ0;�P�<�2Ӌ�x
�xA��֢��L�v���I��L��IV�1#�]�Wn�B0oSGΥH_�E�����*N+`Bq1�b>�p.f�j�c?}�3{Y�Z^@~��u&|���X�s׎(Qm̨�������;��O~x�OKOWkDc�P��j����0���8�?�G_䕱k~��n�WF� U|9�	R��N6m�N��t�1?�6�ڈ/�7:y�c�A��~XP��ܘ8k��G��;e�(��3������N8�:���7�ʙ�9�!G��5~�b��D�j�BU )3�1Vvh�����#���+�+��FۉZ� cU���_tu����*2�$T�os��!��1��9��bx�*j������8^G��5��]�Z�����GY�/�4�\|o���0���1xy�J�������^a}����$�p]'�mZ����+mt�J���d�� �IAc�)�ٰ�����s%���y��a�����G�<_SO�P%fD3��I�?��6Pޭ$|糶�9��H�&���fj7!�_\)�R��;K��࣊c�^��G���z�2n�up�Nd�
v��E�䅧IR'���)��i��ki����N�1W�>���l�%�F�^����Y��M����.�ł⟇�������Q�eSpÈ-�+�{�0�a�)��=����M�	{�RMc#"�2��S^@l�߀��(٣���$��0�i�QV�t���f����wM��M�������<��VU����;1S���^����ha�LsŠ�=���YR�̄��_*�M_7�yӹC�*��X�j?X�AE�4y�3WLt�b_��
�ʟ�I�,���6���K��&�!4'��X�ϧW��vgZ��.r[ϰXD��Jl'su�wa�(�Cr���/2H�k� �P⎉�X|�p\'�Cά?Ys.,�UWP�M�׷ʩ��^�>ǝXʲo���!��J�=:si�>k�"�����;���9��c���Z�wb�i�6$Lq��ԩ��x_���j���R�ԟ��=�>\�m����+� lԋ&� ��^�Q����h㑜}�7�ú R��D6|&]/����%h�_�S�X���X�	ܙ�
��������z�E�G/����lݡa����} ����~~o=f#h�%��C�4�F��>X�#{��[d��+��F���s�8g��nYi�z=["O
��H�!aM`~[~MP�N� �ѲЃF���>^䍂��<i˟O�^N�+�������Q�W)��xT��+	"j�V�]y�{�S�0�i,p�}=ԏ��b��{�c3z��~�qQ?�\�'�r�RE�'�a}t�ǫ���v��|�|F�'��>پz��)MS�.�B/�YƐ�m?�y�qtP�v�P�9��ߝ�A�mI�pm>K��4
�F�OVէ�rL
Ԓ����3��4���X}��ԍ@���	q)?/�. c%u~��{�D@j����v��uT�l�����E�e�lH4�8
@"h��{4A(%	(!�<Nz�[�5MM����/)ɉ �Q�}�,�F��.\�D�]�,1#Y�$i��ۤ��]���яu��K�3Ij���_i^���/�1^�f����@���r8�d�R�����|�ꆙ�2����&k��h�2�"\2ipK��|`,�7�V�1�S��kͳL�j ���"���׳O��_�oh���*g�N
�����B���  ��'R��c��[7,}Xn��إX��d�ޘ2�$m��EzC�.���j���=
jl%(���b*R	�)��&�2zϖ�D�������b�`9(�!�QSl� �j���*#9��=?2���B,��y�t$7Ȕ�=�����{�x(��ϢG2� ��;�|��D��̪�EQ�|
�]�:�$��Z Y�Uк���@�K�6���{ܚO��mv$�S���is��X�@Z��/q�,���߽�@!o̬+:��&~����W��3���3OᚴK��{=���,�XuCer)�u��:���b���[�NLj����܋��ỹ� <�H
��� �W�Y�H��g�����DC��chd*BMi(������T�'J*��k �T��b��#��,�.�7C:���]/ܑ݉ �?P��ٯ�?;�҅���1Y�(��Dp�
ZC��:�c����N�*�b���fE�t�}�=����N�S9�aYV��:�T?ܛ��v`�{�"y�Cdf"j�H�+"<5O�ŖEハ�F�l��i.� ��/s����
u��)�`����ϑ��&�o�,m�O��ں������|�LӠ���:��Uݛ��T�'"x��0D'%���.R2������u��vc�"k���z��)h��w��`�A��  � ���U�fU�J��	�F������9b�����M���W�װ)�+��mr�B�+ �T��/���֝ �E'���t���.\е��6��Sh��̥�=���Ӷq���6.�ai����J)p��St@��ǐh}샀b��^�d"���@���^~���v���a).�U2��
?:����Q<������S},�O3ŮJ�?3�Kb��MH�ؤ+�	���h�!-�l���\w�g�/g8Aף�����걘��K�r�'q��d~d�à��I⎠U���N�^G���eSq�O���n���j�>��_��9Y��G1�}���ǩ�������(xr�K�{8�v�/bِh6���8�V�a����T|\��E�`q���*�F��5|����y`~@����9V�t�����{l�A���   � ���u�j_f���
X.)�-A�uPb�����O�����^�n�Z�h��BU��Tz� ��@��@�dID>ƖM��F�$r|(PW�F{ܝC���?#�A��gt2�-Q4�Or�z�k���󮏞�����}@R�
S��S�|f�5<��������Ñs8����YV�ѣ��;��4��_�q��΄ٗ.'�d�n���(ң��p&L1���g�6�0a� �L2��$b3 ��h̨L���p�žn`ӯ˨����~j�E��"d�B����X��B&?]5���i�e(T��k3%�uw��KJ\�-=p�R����6_��?����t;�y��UL��'�������-i�ɋC3�\�5���`�Em9mc{�e�uM�hX���UDH몘b�B)���돀��=���8��6<�A\��   T �"-���é6�����
&�0�X�Á����?�����P@��ը��=I�)e� f�c�/P}zÔ�� DB���my��x瞠�w������ ���5��>Mm0��V�<	�L����9l'�.��e�K�!��@C�E�ԂV��`.m��3��`/���j�	�wy�H��4K8�F�� r�ӳ� ��=��5�cK���T)
Y.ɇG|r�����#�Si5w��Lk۶��d��<�N3�ࡀ���n��nx�A� ErʷO������=Q{򧪒��@ �M{�(��+HE�#D�Y^9#h;C�	0����_�:����Mq�|Y(�N��   �8����C��Y��1V���ZV����e�o�L�iE�|�nX����F��\Jp�= �_*MQC9��{kIm^2��p���[