�I@�Bi�H�A�Fl�\���}�ђ���`����!��
���p2�;|�J��=��kP_�S"W��	��P��V�tBL��t�.�(�Y�l�K;�Vj��x��#��yێ�_�$M��!Z������Jp'nM쪀%�C�ӂ�Re�KP�Ӻ�˩]��U�/Ґ�eG�Ꭲ���ț�*�?�������ޫ glR��=¥�tΰ!A�5sF�������{�[&.��>Z2T��k��[%L/�A���`1�L��,>\�����'O�7z	��
gOgs�����Ur��tf��	LiDN+!�b��w]so�_���c���1��D#>X�(���w��٭0Q��a��-�F���C��I�^���B��5%D�΀L�,��Y[�v�1��1r�gM��դ����|pd�B�Bd�E$'��"��gg>P��A�;>@��nθ���]��nF`@�p�Ӹ�J)�UL��a��$햣�ϙ~�q�l? �& �U��h�&��5n��^{�j�.�d�RL��w���m��R|�[D��ي?�OP�����lU��P�;�D�2w�����Ql	�":���K�zPܩ���F
���a޻��J٬&��.�b"��9���"2�S�)�hb{7�pa=Ѐe�|�hg�"����=|�L�qXm4�H�R"i���G�Oݣ��S�`�[�)��B�=NQ;j%�6��s\���AYt'�hW˫��܎��T�[�'�K���n��H}�8z�N��.$�|�����F����kW=J�OsuLh��_��Ak۳�3 ~9����S;�iJL�+h{�a.h&�e�L�����$}�����ے咝BLqE��,�׵lO��Lf�T
�)N9��>�Ocu�S�]8e.>�C�v󱥖 ���{#���K\�E�o�v1����\[��'4�B���-�x+����吆����(��(xxm�P=��S[�:����h�8|G��Њ��~�l�<���Hq&��Gi�i�ŋP#(�Ͷ�|�
�B0��S���|�>|d�&��u:��9�UH�����S��Kx�?����h�-K?��;���C�Y����j�3��8c���G|��*�K��c����8�������o�Ʉ��E��@��RaO ���.Z~��~[yfϽ+{�oz�!����F]/]~ !�y�a��͎wD�'2(����� ò�23ـ�IS	��#�.4��RBm7������d���+�5��^��