�2ϰ����(9�PB�!� @��Ja�~8��n�ľ���'�Ps
�Щ�o�GKc�%>ф[�=;p�u$tJ��U���`�崄N��Y�ʛYXI~�IXUӳ�+�I�����9Dȹϒ�"���z����� N�>
Uz̐�H�%1�o���'T��sHL�8 q��:$�رɜ��<Hd�GN�.���oE�M��Hjv3�JY��9(�=|�̿;�}�
|G�
T{�W��g�DH��c�����a����fb���E����m��˧=����o	Ty�h鄗�K�N�;�O���=��E���->á�#-�V�����)�Bn�)��V$�Ѥ�G��]�(_�b;�^	a��� "L�:��m);�%ٮ7X��e0DIדVpTľ:*A���W�`s�$h��mǆ(��Sݱ�酔������A�AUǌ�;x���KG ����]88�f�;�T��')N=��:{�h�}>��^
���Ȗ�}t]*�'U���+�Vք.	�-���E�H��I�;t~3��Ƀ+���=�݋ǋ���̀�k�%0(辗H?V�L��jo���q�^BBR)V��ي��c�{Q�+�����*��ɩ,Q+8~J�e?�*,�J�Ƽ���D���V\4_y7�h&#F!�����lrhZ-��2A}F�`J�sl��8��t�A%�G��s��ij~|�n0��b�3F�!h��)���rw9y�OɨV�mÕ��kq��(�@�aU�[���f�Th[���B���q�.a��s�X��ׇ�Z}��ism�Co[fp���g���Q�Awfd��b�l�a2���,q
���%��\�N2��(���d�;�ؖ������,�aRǲ�!h��:<Ɍ�BXWA����Mc�~a�	t؟] ���$m�(ߣP�
AV�4�x�!��T�>����&�}��и�H�k��&4��k�*Ɇ���n�pY��|�,��(������CEB�6�>��{L�%R��U"��Ph��Q[�d��)��]F�#�aC
�=�,��/��Dƽ��9��Z�B�6=��kS�葁�]��U�&=c��l��*�v�=���xܢN���Q
�	
v��;��'����RI�d��Ph~�ZgA3�fs�з�{�pO�� �,�t���T7Ԯ��)@MƢҟ�j�T� L�1��ԩXcT��\�5�p4�1
mjŕ昲��^&�� ��u�	uv0|}�?]��-�� �h�2���u��_h's^�������Ih'��\��uJ�b�4��^P����,l�_Hm!�=���q���a�}5~�P��ڮ]��<�F���ִ��h�����S����e���~�*<�XDM i	L����}�l��?jF$�ֲ�L��"@< �Xf��_��K=�0H�)��{-P��O�
=���q?-ٳ^���Ԇ���e��P~�>����n4�����o:�}��Q4=�n�����5�}�[B�2�/�ьvg��u(�o2Z�5�*��!4�5
��܍yw�&�׀K�ݲc����g e�/�A����G�:�fz[\��� �_b��QMg.s��V9�kݣ�l1��焯 ��Ž���yVbr�߾�6(��Д3��w�(~��(�'i�����2Ҋ>�tr�c�@k�1�\�������_��ԟ�p%� V5Kx�f�������E5��Ћy9|}t�Z=`��iO�7W�؃���Լ���x(qw_<��Hα�ᖤC~�ib�[�E���4kJ�/��p�p���"��e�Uz,ժ���d���E�+J�t-(yүz�>xs����l�y��a��(��|P�5g>���Uſ�|��z���2Z*S�}P+3Ch��d�vO(��L��"ώ���fԿ��L�l�)������0{��{V��iV��/�O~fi���YGF�] �(*G,z�(!◾��hI/p����{9������fG�5������Y��r�W��Q�e�n3�O�Fv�-uaF7+1�e�'$%{��[Q������m�32���8�/�[q�c��d�N��Ĥ=Ws�����X���S��e�e��xy�:�$5`��b���XIv΍�΋W�R�>��1��g�E\�q�V�h���	��N��|1���g�J�BdcY�8�n�;���P*X*P@��+�����.��d�ӡg|7�oo;��w�ٌF�����i�i�G2.�%Z�iN��T�~b�HQ	��Sx�o|�:+1�f|z��