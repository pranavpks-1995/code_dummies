2�O8�Ѽ�� :��n����v�|��k�e݃_t��U�˲���=��!gB����rs=m�:5��#�GV�>�-%Qw�z��Rd�'c/����hW�U�WNI���+�3��cQJ^�B ^�.����C�]�� Y�-6X�؛�=]q��0�
+�����ub%S�	U�~O��dcEAl#Էpo��(����=�M��~L*]�ާCB)rd.1	7�e�,=��p����D�irk�\��C��h>�`��|�X�r��ns�ĥ�倜�v�TG�ڽ�g�����[�uS��YA�F)� S  !�D�ᎌ,&Y�s��u^&���s,���%tŒFS����O�yXe�@W� �{�A`Io�b�>���s��%�7�Y�ِ���ˍ��
�NP�DU��������D�S;���� ]�Xs
�H/������5��" � -Es� ��C�X�Xݲ�ъ�����8ޓq��o��p�|�]Y��"�]��|�C�j�9�BQ]+e��<�{h�	��ˈ����V)�h�9��Kِ�[њIK�%�[����Q7�7"�Jt���R��4]�=a�*�`� �>���$�C�����p�J{��#L��%� f�N�]��*?$�LE�����	Bt/�0!��񡠋x��N,���߲sB��͟�앀h'�����~k��_6v�H�F�+:�?^g�f�U��P��aH�[t��)r��x�J�Wl�{��D��f#c�గ���?l�@�-&5m���&�BN2�>nJ��?�//��[��2 �'t���絮�9�]����6x�������,��S���"�^����HVb[m�6jO���V��,pf�)�<�� Q�l�5FnT���BW$F��
�QϽ;���ōX?w�f8�KZV9~m�k$�l�ū��5-΄�[��z�=>/�P�3�vw�Bb��BQ���=(�(��ɘ��e��z�J�ؚZ��8���6�5>Q(��'&��+��L�c�Jn��R�҉�1c�>ai�NE�s�	m�	�왐;<��z6�c�^|�����0B����CvѬ*��궠����/A���n>���z��J�f�l�M��p���a��<gW��٫�ԡ����)r�M��b`��-%�<e��.I��j��H�:�= ��(��=���G��[����x&u��s?��\�5X�L5��\��ݧ�z�#�����Ʒ�=�_�QC#��MX]��8������x	��5�-��*s*���BD�di��G��Jy���㡮�3��c��O�9E��p5p7�scmx����!nY�{z
�66��*���v�KB��O/��o@���䮹M-����j@�#'����I)Gf���5kG�T����)ަ(��n� Z(C�T�՚_������©��b��[r�?R�%�1����*ٰ#����nȹ�>MQ#U���z�(��-4�% �#}"�4�L�1=_n6�b�U>ƞ�K�qq�p�g��9�A�R�%���4�G�)P�>��/�d����;��q�V� x���,x�Rh�v-��Eo_�0@��'h�6�7H�
�Ҭ�0�N
h�O��������w��&��uq�IIj�޻Ax.;�֝��T��@f|Aڍ�����\
x�8pT(��{��y��P�>�i�^�KH��~8��L�& j�5�+��F���M&���G���<ڹ '��˳��z��_�6�*�"տ�;���v6&e���R�.���[�UfՑg��9�-ˮ%��� �kj�v�T�R���Yz�ɓh���ͳ�����N����%л[����@���0Xl�C(z�/ʣD4� *  , �$��,t`����%Hh� ���7m��x����R�YYy��ǩ~������ ��;m�����G��'0��E�c�������y#��j��2����&☘��3�S��$*�g��=��9O��~�1����wJD6�L�-濍遲�'��F��񡪋N�����v�~e�Z�@��X�ރ���w1V��(9����0�4(��,�;A��&�k����ޫy��"���a��o����?ե̎�]��%µ���'�5�+���#h��A��y��t��7�=_��[\���6�,�{�x���Kֶ�8�C�Ӡ�SYg�+r��m���Z&>uЋ���|AJ� TJU �}=�hU�GZ��h�Z����&8�S����������LKC�t��D����sY�Z~��ɀp
��-��1X��{�|�0��4bz���j��K�N8N�GQ؏��1��Y�H<$��5Px#g�
v�`F��~Ɵ�;3�W�||��&	�ʅ݆�(���T��F��l�=�ٽ��fZ�"n�3N3��������G�$��ۈ�0d t&Be��|Z�{�mS�5�&����T���Z��7�5����<�M��}0��/q'�w�~;G����l��	�%�t�b�=h�S�6�ƴ�6yD$���������>���~�k>�v�N��djc=a�نF�ְ����P���fMhA5��'=��K�/B	�0�
�Fȹ�7�m������L���0�� %r�$�@�r\7�ݍ�a���붩�)��aJGZ'٪��T�F�e���^( ��s,E�Aj�>}���.>F��²��6_��0A�<Rxǵ��Sy�N��%.�,wp�Q���ձ+M���\J؅>s~l�:xD���TDj�~��4E��|b�W�W�s��-\R��p�NS�e�WУt7;8�/�e��z(�-=�-g��Uҫ�;�(x�69?��B���CY:7S�f<şA~;*Y�  ���xU�&�&+.6ٝ�k�����]1��|�-�5��W��p�_́N   ��@����c���� �;A)Yn��⢠�GNe�ɵ�\�T��a�yI���WP�p�H�z͡��8��0��=�9]-ل˃�sh1r�-+<cs��c�2㺲����+����J1�v\��-B% ���,��xX;�{��;	%<�m�����D��8�m?4_���w(˓�Ŧyp����&�C�L�7�\��f�5�S�-�V��h�~˙�3��t|O�d˓� �1����Eݼ����ƚ�D�c��A�7�2Qe�B�6�d���<��� 5Pp�K��if?'��[��iN_Xk�:��K����̂����>z�l|:�cU�o�E�����2�<ҏ}$�<�갢h���[Q�=��}^��SN�Y�f��ǐ	�x�L��+�Ȥ;С^Ks��v���.\&�)���ǹȺ�������E��zƏ��,���Fˀ�432���*��O=����Ӊ9��Q�i���Cn�RJ��s�f��S�0�>���~�������~"� ��������JG'���V7��W��,�r�-Y���i�$c�a:�`ҽl*����rB�'FƓ��G>�)%��	I�x�"�2/��Lv�r��y��v���G����I�Ḫ����^+���NYS�q�:qJ>� c�����נ�|�n$(�(�͒����R���&��4Ŕ�0��𚐏h�k2�t���F��m!�fA�h�#ȫ#g-C���L�>�ʍ��^y�<�in�����Xpn�f�s"&��ߡ=K�[T�HEc�c�DQ�9h{p���G�2x6"!ג�k��hD��b���*����J��#�p�^��&Dg��#,�OG,c&�f�%���_RE��_�B
�=���d&�J�(ׯX[���=C���2jL�0-�d�	���EǮ��BxY���/�)�堸�w/�����v���u��nC4�7�|�Ty�Fp�'FܣmI�p�xi�^���ks����=�6��!�3`�
��Nh�%{�0�:Q���Z�M�7��.8��f��}vj�ˊ���6c��~)��̈�� kl�H�����UХ}S�jA6��	L*�(so��};<������R�fz����tBJ��|�l�h�^��������^�d�J���t{��~BɨW�/��,ڎ��������h�+e�kAm�nJ�F��d����e�H�u�sl.���){�"퉠����'>X�\�^?�^�\<�ek=r�j�%f?���fWZ�E�Pr��2��	RS�^��ч-^H(����#�`XJ��-��y���֝�̝�X��!p�^V��t����.3�!0�Xn�ri?P�H��785^ssV*WIp������E�T,��0���=�5�$^`t�R|���]\-��l ��� :D�V(��E�`�WS��U�┯�1����4F�����O���^���O~d����ǔ����n�!�&��h���F2%"haA�����0vʡ��A�D���M$��L�����@���R�L�����I@�<�L��_(�o�T��
��:�g���5\\ҟ��q~�|��[��,;.����{ge�JV&��a�hb(�LO�K.%�KM�6i�mЕ�Qa��d��x�-�#ulc�$u��J���֐�� �,�cV@C�B�|�G\G�Eh��I��BE����O�%WN�0��~
9_gO�8�t��x�Q�>[�s���t�R�aVp���"��>$MO�O��@$���ІŦL�]�7��3o�ڏ�C�]�������yJ;%���|%�C��ci5���|y�l���W�LD�㹏w� 7��[<q�q�!!�����(��d*xR��C0����G�9M���Ӻ�li�S�����+�D8l�� �`�0O�í�CuB%uF�іh10��]v+w�	�����d��s���� B<Q�����&酟Ҡh"�3��=�9w��(�ъ� ��Z��[oic��^}��`{�Խ ���z���FI���q���
��_RF�k'3sJ�bb@�WTy�Z���d1��@Svw�t�����n{(�XOg