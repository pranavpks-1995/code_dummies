gjQmC+�N�2�m�>�q��x������烯������1˓'-������TB�9�N�Jo</�,nΎ~���髃H����>���"˭LA�GR�R�5mR�M	�;�a|�o����y���Y��g�hY�	00��8c��A��G��-HF;K��-p0F0��w�;��&�\	+�4�$-%��^p+]3�(gZ+���2�s�Y/��R�':C6��ً��N7���BW�Ԗ�C��q�YĎњ��}�ᣍ����o"��T��֬)�S� ���PT�v�]���������I�h�&K'�����W7W���y�RznJf�1F�g�x���2�m�J�3X
Y��ϭb�)�Fsg|�/��W�.��)���h]ѳ&}���y2�&ZP�	Rk�ҭ�E�Eh�+[ԟ�/T�m�-%W}��Ł}{m�Bw�w�~ v����\JWý�Q�N���qc�n4��z ��&�}o)+&~WJ���X�G*B�3Р���Xy�B��=\�!�S�Bw������љI������w�"̏�m/M�h�Sf��yFk���#*"�47�6���o��Cܜk�v]|�n���܂��nV�9���%�O���P����oË�07�Av� *  n ��_��F_������6rN0s��l`�*�.����(��P�� �9d�I�X�/�K����~�v���X���)�f�jQc�i�}e��s��2Ľ��*t�A6Cj�����]6;-� u6qG֬��)j+���V7!�o-){�>4Vp;�nܷ�(���_���=x�@=�*x�����4�]�u9� ���U���5������y���jOhu#���s�]D�|	vnU^�0gd�8l�$nǅ<�{ԩ�}�-Ẹ�݄�����E�5a��9�K�2�t��g�عޖ�!��+VP��g�i�����:%)ol�3��'�k!��&�y�·��b��-@>-�Of`�A� T   � ���_��F���Pf�	�p�y��[E5��P��{j.����z�h������Y������;������C�@��H͵,�΀�Ps`i֑�!w���� uMJ�K��b����o��r998��r���뺞1�&Z��Zu��Q��ы2�1�� {3O��3�
w�5�3���Io/��aS��m�O��;��!ܴ����.<�!�'�S�Epɠ�,�牳G��Gk�������x��cH6@7�\��X��9�3��!��N	I�60kF�+�����ӂv�s�f�ƖO1�������ӓ�*�o>�=���f�5�t�dШh�k`ŧ��#�nu�sp�JR�^e0�N������D)H.o�Q��c8FHC��z�a��8����?�c\�m��Nݪ x(K���J%	l�a�;����؁JaO9��v��ؤ3A)��w2���k��l��-� *��2�E��[@�vh��+Js�G���|dd��տb��B�� �   � ���F:0@8Pں;]�P�T��N�OZF�"r_�.cfM�"|l+�؄O�ش/�s��J���G��r�pw��(�gm��B�*����2�m�AV*�c�t�`���q��.��4�,
![�����\0k5Z�3/X�H�Eg	�O�W�Ԙz� Nd�tm��5�/9B���Z��`��19��y�Nث6\��$���.�R���7ZC�un����SX���s�m���������6��70�if�'`3H�,B�=	���z��0[Zh�%�ui��E&��	�w�rfx#+��\Y�����M\p��*�pL	�=捡S��a�m���o�멼��	�����]Qt�p�[O�ue�OXK�<q�y�%_[�~�#�	��j �yE8��C:!}���/�Ժ���
y�G��i����c)�0T��qs�8K[�?�a��U1n�@:����'�HU�W���-�;�0