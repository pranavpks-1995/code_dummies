!�z�3(�K�*iwH�..{�ZY^}=��mQ9Qg"��Լ�,r{���:�A����|Oa��ȅ�Y�W���&1$H��e-}�}:�QNb]{'���$C�XTl#��5�׆5v�8���\�n�)�����ج�牯!�&�&�<�q��rd���yX	�����G�]V��v��h�`���m�a0�t�<�߳�Q�i3��	��ʯ��+*��ED��r�z����u�E+�D���/s�K=7ߡj2։�~�v�=\l^���Wm����g�=폀��q���X���'T2绝�{��$�:AH�0�1�'E���|J	wغ�@:5�=� ��F�c\��?p�7a�Z�۞��㍔�
���d�6�J����M9�a�͌0���j�?��T_�W�n��ީ
�L-,��=�S0�p�3Ѯ� ӟ�[���YEP6>��r[u\L���/�sޣf-��Zz�+U�[��p�^�����D�፶-��F�pu� �K��^�9�rO��M�ՙb���J<�+,��u~S��T�.�f`� ���ڗ����s�K5	y��vqY/�4�:��H���;�8�?z���_F����zn���Qr��^������n��P����A��ʉDQ5;Ozɣ
�635���f��C˒��ª��?����:߀��X��a��ݏzvґ�b�C���}u�K��U#�;��� ߀�P�=�C �y��nھk6��eej׸!���|�r��0DwrZ�hchl1�#��1H�lA��9�啗w#��[_���r�>�1΀H�����rZ/C_��ˌs�d��G(�8���k�҆�-+�4i�[Bd��wZ����w;���*%�yHG�3�2s\��2������h����#��#9bm��$2�l7�6;��bF�:��Szr�9F�L##A�S��ҫ�-�AP�ߝ1�L���bZ�l��ٗs41C|�*%�O�oy3������pfY����K�.��k��7Q��MLn"��g@eK��<�q;�x�0��	R,p�����Ї�8z�xſEA��%!�l�_�I�q3�Q:�eW��}D�4�yѩ�1�r����m���/�y˞Zyu�X�Z�[��*=D��Tb7�U�"���ë�a���v?�+"]�i��zꀺS�6]=ۿ����z{AM�W�Z6@IlA]!��3m�8� x�Agr �z����$Fv)z�3�gB��4�:�Z�E��d��2���>;3�,T�W%�I�j�