	��w����Y�r�]�v���ڈ&��=F� nk!���aρy'*Z<��!�> ��Ή�,h��,)�b��Y!n�5� �ߏf�TP�T��v�ɴf��C$�
5�A�"�H1o���:�Z�S'ƺ�����Vu�����ɛ��$���*�T|���e`O)��y���=�|0��|����ܾ����x]ϲ r:.�j�[W�`Tc��d��9�V���ƌ�I;)ع�З&M{&�v�[�� Q��J_�G5A8��	�l�@՝��7!P:b�Z��BUw#"8��B�,� ��w��;��5��U�4���H'�����ָ١Q�y���-�B����	F:�Uh	��E����1AD~@�զ �a���<z�T���U1Hh�A罉ܟ�����G�>���;��;�o�,3Y�_8nT�;R����]g�B!`AR�0ws��=gDft�� ��}Bp���V�<�fZ����%3�t���ƷTf5��o��B޳ 1�6��[��e%�ܪ�0��kG�+O-x�F�8*��}�;s�9���4w*��6@���ѫ=�
ג��e�P&�w�/q�M2��Z����I9���# �I���[זv_<[�n���~�spD��#|'����T��� td�Bwښ&܄�B?T�t<nWB��bm@�甡SZAݺ���j�fݷ=bP#>���,�7Dn�ӘYz�֙A�y��i��1��^pcfwc�'0��_V����aEtY���pA����D[j�fW��V�)�!niNx�n�Ќ:�!D�H�Q���F�r�V
� 4�4V.pG:�V|Rl#�:���D�����dhÀ-_H;Cw���|p	^�(�"��H�#�%9E�pN �~��5l�6"�d>��D�AP��>�6�l3��Q݊A���{��{�P�K�8��L����p���nyGfn��&7s��
����F���z=/D���2̧��t%�Xu��ˑ�!J��(28	��2�x<%3��t8�#�(8�M'��u|	���!e�'�ae�Sfl�ݯ��#�&�O8���K�z��CM��0P~}�/���`�7��8���6�\��]G�Hú�_~z��K�`+:�ګ
�o7�6�5�T31��.��$:QBý_񮌮=�9���>JѬ6��q�~r��tM�hȊ07|S4���1"���i`�{��v��㖦������)���Q&<;�;��O=����0�a������K�j�d�M�(2�WatT���E+u7\��)�x�|^���[� �@4