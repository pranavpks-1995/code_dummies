My������r�d�����?��+w���e� 	
R�*�U�ٞ%�"�"�E w�9|d�#:�!�.^�:Ӌ2�es�ӎHX� yNMlg����՛��6����*�+0��^�vPz}�a���N*��P	���g�L���vsD�>'�gVobgguȯ5�|'�OcՂK�S'!tK�##<���S�tQ-�w2�~M�Q ��7[W{nDpK7
)���G��t�3�ՁF:/�1
k4�K�D���ڌ( ���&�u�d�b�h�Q�����j���V�����J�ڟ�Й�Z�ì��>ZaY� L��݆�b�GO��i��!H)u�Kp�O�ZC�k	��[P,��U���W��Q2�/�e�<6��c巸[1�F��-��}��Z�*g2 h��  �+R�^T����ܨ�
)R�?�֢�Zm�Y�Rc� l�<�Z�P��it-j�Dp��l�d�lζ)X�D.}�t"�#�-Z!�غA�����Ņ�<����U��ꤦ�a�-�����>܁�/!�F����]�^��v�Cn��ou
��F,��Q��p�jsz'�w>�����ӏ�����D%"H^���vA2�+i���K�W;�|�3h�s�l	{42�*�M�R����c���%*�/���fՅ	g�.iR�W�������Kz�2���e�l����?�S��(������ iB%�/�Y����n�u���FI*7K��͜�9R������?ӛ����Pz�-/n�U?�=��ǐ˶Z���ah���dG(n�(�\el�NHS�j�z���5W�E(Z>O��ᕛ��������
?TwlJ���w�,�� ���<
�J�u$��,[%#̝��Oȸ�E�^�L�}�f �'��雹�A/�1%`@>/yAh�� [>��Y���͸�z5�3�B������lx��1bЇnT�j����nD�7�`��
|&o�"�r�!�Q}�Y��l��nY8��4�����L|o�g��6���:�Q�o�w�~�b�&XTf1�"�k�q	�)���.�����3@dc�ʺ����j؂*i�l�jp9��:��&Ik�Ek�:��}�� \$����B{Ϭ<�UEL!̼Y�3�j��ܤ�u5��'{��G�&�l`�Doڠ�6������
𶱘��\m�z�,�o=|W4|v<��m���qN%�[e7�ʤ�����������ߟ.9�=�@�*�R�P�Q+��2���x��DA��w�#e����zh,򸮱}�1(t��6�+�9=l��}��_�@
Eӕ�X��N�؞+wC����}jmR����o%�k�e�
�D$�
({!;�]I:�oI�T�6��
)�Q��Q5�z��aܒ�P��]����iO(<5�dL.�q�n�r�