c-�۝�9�r�#��~<y��*�����v�.I$7���B���ج�pʏ��-]J�k�èc����S&2}���6�4��YH
-)�5N�̗�SS��:���.>���'�]�íC0��(���8����NV�����6���|���A����F@��	��9S�R�Q&Q~NJYLC��@�l���^�Θ��^U�_����Nçca#&�|��}����k,\��W�]:ԍ�QD��3q\�i�ӯ�f�bv�h��ͱ@����C?�4�����C�0��VqU5�)�7j�	�]%0!�!v������M����>H�i`�O���@P?�V�qO�̵��$�N��������S�g�
0U���t�� Z5Er����4cf���c2KFC0��0����" |0'���l����`�(Tk2zӸ��i���|��[�}�e��N
*}Z� �꽜�	�=�v��oW�Y� �����u"夠���}.U<����t��l�X��*{��p���_Hz�K�QǱ��&�h|Z��$�ƮB]��3a������v:������~f���bJϑ}:Ԋ�kGȭ���ʂ'�Ғ�����c����� �6�"�}�?Q��(U�Z89�(���_�Mu��"���=!��g�=�cJ�NۧJO��<�@"�I�~�8o�0�5������S��V�}���46�L�;�T/���\\�%��Y]��[�X�����g-1��m�<7�t�ّ�g��];�j$�g@�p�bW�����
����a��R�M���?1�}):F��(�_%c^�P����Ö��k�]�gV�t~p�P���F��9t�eA}u��v_ 0X��͉+��J�Ț���JФ9���������8�����Kϟ ��@�J�R���;�>��xj�����x���ƨ���	ԩY�th�	���7@�����%��[W8I2ͧT�ߋq����*�k��� �.��_݌d;����;~'9qhQ�x�v#V�5{�j�p�d�GM^G6�ݿ�<߁�&=}�@�E܁  � �f���,t`���9�Tٻ[+��m�<��ԩ|_xn�'�Ƹ�=Ѻ0qZ�樁�E�f�:�XWzl��o�$t��?�ܶ�Q�JU�ɟ$D^��paT+@9�& �'F�}�Q��k3L��>v��-�!���bB���of�d��ČE�X�mJd�S�⬧�z�j�z'�D�FYX!�xB��<�L̍���X���Mi7��(�g3c�;�_�5�#��p+g(�Z�cQ������$�T����&p:��$mb��{�o�_ ��U��M��tJ�����$h�2H�W�v�(����u�ջ_I�4Ov��>ԫ$����TUe��Vف�N�)%�v�����h
]me6A�ⳮH�YeBS-�"l�듃ۮŏ�s�����w���X�±
8��`��s%���`0� 	�/U>�.�MŦjM�t�m��1�l���u1H�r�C{��?����l��>�M"���\c��#�	
C��4 @W�L�*��(� ʔE��� F��DMkU�YF�Ʃ���lB����O���!g멡��(f�Ɛ�]���RB.Z�F��? %� �+9����Z	P[S����@�z�dV�:�/���2)lcl��u8��O\�S�VU��+��&��vC���"X�?&>�����k�~�:8s/ɼ���0.�$�ܾ�
��7��t�r׊^�zd�{Z�Rз`��P`�\[Y��)�Y�.MP�r���/�n����̈ꡃ&`ŖF��N�]��QDO���7f�G� ��&	��#&B;}���~�>�eJg��'�ěQG�.����������^c[���o�-����60�-ک	0�3y�_<�D�ۀ����_l�$<�G[qA�j���{�;(�{D�W�3L =�/�F1���Sެ��,���Q%T3�<�z��������=ȡ�$��1��F1������/"ٱ��������ǀP/.�Ph�^%�]�c���w ��^�E�e��:%M�	�A8��|��l.ݡu��r��Dּ &�qF
s0�×F_4��ӳc�KgL�_���b@|�)}10$yE���O>kV��I��Ő�������F�����J�h%O-l2o��r�ė̳2;q�� ��!3$G��'����_)�H�U�Z���})�k?$�^T�w �i��@j~&I�YLQ�����r~F��?�`��?qs	Pf���I:�����������K<��<��8�&K��鿑&��~��qgP:�)daZUsj�}L�a6����܄���_L`��z�C�o�}t��zJƆ��(��];檐̈́,�#9��M��8]�U��~+*W͘��$:�
�Bh��Kt?����0��|��$t��=������QRLݎ!�}B��[��}x+-!䉝�:iO�G����)�.a��>7O+k�uM2�-lh��`E������(%#Z��Yc��o�5mǂ��`e�P��F���Eg�o   _ �-W�������m��v�'@6�Q-��Ϙ ���P��s2j��P���x�)�]z/CrL�QŸ6C+���Jj[��4���4 |���?�e7]�=m-�2Qˬ���ou�5�� � !�L�zY�.S� ��Fc5o�w�� ۝W)FĜ�_�!�z��*�C>����C�"EXd��_��V̈́3=�Ӷ���a�>p(�F�3m͓l�dj9�55�/�[Ͱ�]�i�@IF��#������9���Io�-0���ܧ��� ��;�%�K�<�)]��|�"55e ��/S���x����L$Ӭh,�B̀t�1HvUWs�6ˍr�t;5Jі)��ױ��y�T[J63�.A�*�;��GX��
jחN��[��7n-j$K�1�T��#�1�#�nk�2L��d!(x�JJ�P��"NoE�
�KL5ͪ����q�8���F�`�0n��v!��|3�z����jn�M���]�WSӳ���ZѰ���U��3� f��[�%���tY,l�'���!1�M6�퇔{������uA66����b"����d1y�*c]���ä�u�;��a����L�=7�7���y>[M��*]��12��r�×Us�+�t��JDҼa"���i�*����/)�h��}�� +�dwgH����U�y�J������y��ae�t�R0�1O���ܽ�0s7��׎a��3 S�o���= Dn���� <�w��5�>ߤ՞8*1�Vm�hTjjE|.x�(�:��5j	�ڶN"�dBG�H�<si*���������n���ٍgV:~h} �ΆV�nr��.[o���5�I��-3�O�{u/nuM�T5��x���d���y�^]�<��BW@��5�[&�Z �e��!DhTPڐn&Q�=� T�0<BK��(s�����!h��@wN�bL�����M�̐#�;�q�Xq�H#t���*�D�r��qN��a?L���w��`��l<H6$J�@V�����xn�|-�������WK�5W��f�H�����3k�z�����1��.xx�v��2y�w���#^Aby�N����庣�ZJ�"�,&�N����?�bՕ���G
�;��z�
9���U*S���8�6�B�3���%e9O����G�:w��F7��0(��P/��+����A�6�3����v�XDb2�~�y���9��J��ꧽ�OX���<6t���{_L��T3��{v,�'X��j����0;!�A	5�� �m��<��s!��k �Jf�"�4,�9)_^i�����P~�˧e�h�g��dG�~���$�娀��4�E�d��Eh������Ǡ��!��$���";
��c  Z�s�kF\}�:���&?S����V$:eXjqrw]�Q�̤e���� 5������.��u������^��v�$kZ�aap0��{�O�A������th��OT! O�M�[�I��o���wr:������     0 !��Ƅ���*;	���lҬ�MU�E (�rN������f�M�=�h�0�u�.~�c���(�T� +�keb������#9~kx�dV<]��*>Ww ��s������d �1��	/����*k]__����Q�pտ�Зp�P����7�i�?y�G����gV0�    p!���C�L�T�f��P�a}�� ͒�6�<��4E�iF(�θ��-�:��c=��í?Go~+l��(�q�r�Ȩ�i<d� �P�/��&��ժ��%3���k��쀰&ά����$��>����	�(|CT/�Y5��iW{y����7n��     p!��"š���ao	`̺���1hU���O��TTp��B��Q�[;�=�`��a�]����m�> �O<X�����~��on�W��}t�5Y�d�>Uc`M�� q�&d�`�(�٧$�l�k*�΍7M#Y!��޾���H�gtܢb��	��M�N	C�e����:�[~e��qv��-��?s�     !��.��D�l2*�^A�y����u���'�h�-�7>�,�K
z��a���m��ף����t��Rb��!���� X:�1�hCiNP���e=J��_���B�����)-T�-�c�*�E@%��DtR �<{����+ֶ������0    8!��!��0�a���⋈�0c�ܶ�|���\ږ��@�I�)pߥ�qy�\9��27;�}�'qۭ��\6������!9_���u�|�)^�=t����ۗ�.�m�D;+����r��Ժ ��@
�h '�a�[Kw��D�O�cT  ��!���ı �Fr$�%w���(E��=������2��%sQ�$�s��`��T凎e���T��kz�J�� %�\��4e�vfd_�y���K&U=GYg0���8�&���L��hB���  �N��<ޚ�`��B}y�bS���b������gѶq�j��    �!���±* DW�  �,o&.XZWR�9�`�+>.
 sU���h��>�������s�������:h�����80K,6}��c���˪����_��*�$�y?���/���wO� �=?�0 �� 	�(&�B:x��~�G�`�x��'�u�߯4��� ��Rȁ@   ��вUW�C����u5yo[��V`�=��&�+r���F_z��ܔ�StF�a� s�?�]q�>�g���m)i��ZݻK����(s�:�@�IH�F�[�{vr���s���;�me�L���:��F03da�����ġ���m�������yÑ�f
"��m�]u9jD�N�Jٸu̠��<�ﱓ1`d����_�r��y�+��K��R�c��߆e8�?#���g0`�����������/rJ����$��Ы)���݋8��K+Q$�%.Q�.ܝ����WJ-����gD2�m��;i6��O������dB�4X��O2Ǎ\��Ϸ�	qg���_!�6�ϑ��53^�)��'��; uD�Iˎ���|����Rg��]zL{����4�[WD�&�K�ľ���L����*Wr0��l�({�2���KӐ��i�:s��Z���v$;��7%����h(j�� w~c)t?�]� ����뾓�R����'6j�3�<�/O�_l��V6=x���"���Ieh��!����`J<X��J�\XL�Ҫ��YN"Y�q%��ȕʷ߲k2}�ʝ�KRxoX�3y}F���+
O�̷k�
?��(Ѡ�(HRU~p9���s;�5�}]%:��uph�zg]���?�v��p�?�&z��O�J�_��#��tYj��"ҮfuEƧ����%7��RP_��E}���U�V��ݺJ�����|��9�4���_[�f������y�f&à6c�E����J}r*{�b�����D@s�R�������S;�2�F�@{a8�UJ:%����f���#��E4&��W�rb�Q`jO����JXH��|�l��KtG�Y�%������0���g�u�"��i��w��?!+67_Z4���xkp��_$�=���Q궊�i9�P��=��rV�0�_SnZ�h	�ٖ+4�gS�	�� ��Z� S��>8��&~/�21C��/�&Z��\�Q��^��Tm�Z�G��gK�')r��/b�z��ckF�e�*)�0�{�]I���O5�5eQ�M� �whZ��� �ێŉ5��Ǡ�����hz�w�c��c��a<I�<1B��9\b��ri���]�΃3 ��ΰI�����H��R3O�c�\E��"�[� ލX��[�n!�9�=�㬤�?�'�y��+��Dg5T�\��O�Vx��?C1w&�p]
��54��E�^< ��ϸ��al��v����M�����#7u9X�|:g���"���p���Q��-��n��T'��^²�.���B􂺗�_��[�����#WEr������X%��L��b�����7�9쁞`C\����Q/@��ܴuei�MS��u�'\���A2������\>b҅�BK��^ą�AIDq�V�.�,����pw�����LY	2�i��T���l�i?�C�y�K%����d�(Q���m�� ��|cѵ�x�s�	U�,�F����-é�4wU����0|&��˦�L��NY��̄�K6*���"ˈ��k-��G�S��X��.Ѭ�a��� �Q#nQמ��X���OQ&��ӆ�P$ɩ:����yF|�Ta��dU[���w���Z��0�\>r����E`�J|��>p`��:��E%J1ff�t���n�e���l�뾴R�>����,��Y�ظ�i��'�Lhew�	��3Mt�ˢ
�ě�W{�`˳]�:'_W��ȴq
8W��Xq"-tӡC��4�/�m�P�^��5MK��2(��_�5fa��m��1�Vv8�q@9	�� Y�7��?��ǔ�x�X=,�D���]c��u����4�a���
W���V��j�C��_� ]pŠ�Y&۵���ɳ�����Z�����c�>���L)s@F�y��h>��XZD}w�s���E=Ѭ8�+*�6UB@KYZX4�����xob��(ܔ^=�)��������� _����]�<����B�|%A���RY:�������O���n��w�]������#��a]��y��㩝`L��(��nC��	܌�1r�<�-HБ�� ���mx>PZ�<�as�I�`�4�gnh�0c%�o��+;e���������x�@v�4�}��B !z"#fGX�p'x�m��ł��M^���W'�r �ʁQ*�'ћ�t����u��py���Iq�e���;
�+�Z��N|�1�w؞*M�7T��і������v˲V��ĶU�|�xz;�0��ҫR۵����U5�*&��&:-}s��C���K?%͛�����w��):�g���1�O�04R�4Ė�#�s�ػT��N=�bA	�凌�J�[f�z�*/�yG~^HB��?�,�2f��dD7��g�4�+s����q.bi�[n�iCN	�vw[��(����0��y��dZ	h��[��!t6����IGP� �=�Ν�;+@e��7�eS�L=ꊅ,�b'a}��Vh�?�@ �ј����Y�.1�ت�;�_��#����0������>���W7<�4�A����`�g-�D8p_�p�t�үc�vr�]�A7���	��֫c+W�?��M
5�0Vu�pBNӻ���o���s?����������@p� �	]� �ȡ����(�� (X�s�xk
P�Vp���Ɋ}hʇ^�Y���(�n�Gu�F~�[�~i�%�Z2�ۡ�ġ��I͔�\S��z����{��9_N/���!Ϥ">�R��>�i���<��A˥���a%kW�$ǙD>��	���1ʓ?In_�^�&cP\�N҆dR��@NQ������z!�+ݫ����g��C���b���/�Kiɡ��Xt��g���N�0�F�C��{�ߴ��Ÿ7ҩ��5�kN�j�X1�i�Z��Jz|��fGoK�K>关`e��G볟k]��>�msP��oʨ칙�֚Kj1L��7�_oB"���)�[��W-�yv��e����˓i~��U<?H�����13�7����$oY�">xc�#�	��X>ȻȅMK� W��V��z^��3y�"|����!�P������X�SU��^�a��M������F�O����&�@���\���0
����'Z:}"�L@���W���}�y~uh�|�_���y�JS��q1Oj�W=���_�c�6��t�Ou����G@��m]����8vt&Y�j 1�t���SU	��y���ʀ��Bn��uY9�l+��^:��s�$���}惬|���@��{���
��u��^r���I��i��+�-G����ǲ�k�]�x������؊�ER28#Ob_�]�Z�;���U}�a}�t� �q�8�D��t�/�q`����Ĉ5a�Z���"˾�n��vQǵl���>&��0Eacs3�+��'�eW������_���~�x�(���Z�S�N溃� 7 ��ˬ�w&��Cr[��ї5���tO��g��?`��<�B��ѲA�)��g����IU\�5�͔]��ŏh�5��iË���d*�ؔ��!��g"��\6)U�
��}��!�����Gbs���a���&F��D�d�]jF���j|x	�d��y0&�񰶚6
�<&��`��U��V�c�6x׻DB����:��a� ױ������z�0�"U]�-L��9��&�������3`n���T���1a���!{�A�����{�t�N���D 9��l�c�Bq6�(�x��N�n����;y�oE�܎��|٭e��]�pr����������ǝ����&��OK Vw����I�2&� @�?%�a,�����s�1}$s1�&�xq��Ib޳Ɠ�_����T^:/��v�0;� Vr�u#����U��1E�Y�g�"@s�A�#�AaȢ����j~���B|��܃or���?�� ���WK��������f<��|���)�#�::�������e���[EݐʁD�υ���{L��
Mē�'����g�\���:hS&�����>�ruLyJ�]K�-���\7]��{S.��ls�>'vSL��@��_�5хU	��Tİ'7�"(���y|U��Aoq�nqa`&ڑ��:5Y���T8(��*D��0# �bc쑛z��w�e����M�9Ե��T:����b	=q���ʘ�M�3�-�K󒲡-4�& �E+�v�hÁ�C�� ��͠��"���aA�^�%4� ���KjF�7l��I��~Q�=�ؼ����į��cD&�Qw���W<:9.�<ɵ�*�z�LJT�c��J��w���Q-�D�����,� X�06֭Y$#6�I}�P��u��7eg��.��T�ERW���%.�pS5.�l5R��݆����cq�*�~�S9�e>dQBeKx"�q�ܳz9��5&��98\D8�bt��ۄk$7���z�W���A0C�'�yv),�q��8(𺔠ə�-�sS"X?����4p�Dވf0V�Ow�����K�v�E�hj��|/&���F)p���2������"���v�H��T-�d���$&��䤙�5�1sE������7t�Q���&ӅHɎu�ƫO�����4�1⑖<2G ���2$J{x�.7��G��蟻�h�ژ��<�~�Q�,@�)E��f����R��&N���OY[W�d@1C���G���  |�%RW�c�*G��Sk��GO��T[�n�MTFgi|��|7� ���[��,y�Ȼ�K�<,���A��:[��ʌoD2r��K�pO�Q'���ׅ��W��߫����

�hչb\(��\�_�ѝ�t4��bo-�k�<A��	a	F�>�U�?KCњ��tǫ!��#�����&�b���8jt��ٷ7� �\�u�{�î���gf��iF�P��n���f���N���x6��c��u�w��,USK��'v�i�kcτ/�f#=�դ�Y��ۓ`4íe3����Vw��?�� �<Ň���O����nN.i��˨�����!��O�I�/L�~�4-��P����G�<^��|;���8|���(�:)��shf�\�7l��~�پ�
v�e+� ��|������y������|P+n���²!	ư����t�l��SM����Pl0��e������2je���3���=N xD�Q
���=E��qi&Я1�Ig�� a����Ap�J-w�>DZ ���7f��Ɏ�o�M(���(Ȕ��&��W�0�����#V����^
�-2`��oc���p�}� 8e�3�]����U����2q���S㎕��ľ�\/�a��H���n��:-(�H�%|� ��N�yļ#E)��HF%�F�nt+sh�/�}���6��݂u�Շ����{zˈ6
�'3�҆���	Q��2+ϕ!�l�!z*��ң�V��}&��ۤ��x���B�5^o
�?K�9ˎ�4��a&1A�g��-�-y��Ͳ�
%b\�柖/ex����5����AX�D%%ehѱ���cN�B