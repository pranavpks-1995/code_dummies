��ԭ�%�^�a�r��c���T��ں3�������ڛҙӷv$9�5�F��Y���{|Թ{\JSI~%�1�	|<�B���l|]�Y�f&Y����[���T�S��@� �j��=��!g��v��ˆ�#�:��m�!W5LhU%��q��V[-

�"z������R�KI�ܰL�"�5���N7~��	]�a�:%�m$��Q=����^����d!����٠3D�{3�-�@u{��dF˷`x���_ӯO��Ok��I�_=v����JE� `�7"��أf��ٮ?t��[���j��ҘQ^#�	�B7����n}��)^��PѺ2���g� �������ın�U���g�p�6Pv>�<�&Qc����dzv`���o[Y��<L�h��"��J��~Z�k�� �2���ᴗ�E����g���j#[y�&��j���՞�L���W���D}�\�q�<��^rb�xFO�����>�=g�8S�q��/s�Kx�S4ju`���w���m���@O�?����V��X�#/)_;D�=~8H\�u�g(��������.��+Y�g�E�=]B�>c弽�W�dI��2̪7��F�u��߉�+�cW6��b=֚5{�f�5�m�CW߁�W��ظ�h��K5;���Y�����P!O�qY�������4��J��r�J�~9�-3CS���&��Ɂ�e �,�n����Bݤ���V�����+���@%Ei���5�	AQ �������g܃�E%{M���k0s��Jg��[/���� @ȅҬ5y��l���	]guo/_z��I���8t�F���@�݆�ŤȮ-��ϛj���^2V��|h�'�&Eʬ/g
Iq�^�\Jd%Sk�%A�|@��wЇ���5�}'c�N7���Rސ����`C�<��"`kf�|����L���!����Z�=FxZ�)�y?�kR|�NH-�1��fJ���r�q�{��t�hK�cd^����-����,�?�y$X�Y)�`{�K]e��a���2
�P\�^���-���-���<<0ɳ�-�RT�/���2u�����}���ݬS
��oj#dd&�� �V`;��E�h���kՋ��g臰4v��_|�5ǳJ+�l%7|?а�X�����crB��4�Z�*�5�NXr)j�#kVv��B
��wqy�|��8RD���Iw/Ǖ�\%�#���������iS�`��y�];�\-y�g"!�3��	ߍ>;@*��NxK}�~R��]ġԚ`�����ő�֕��IO�{�>s
?ol�� �������R�z�\o����+WP	o���J�}��S����r�~����(z�@g[����O;q_( �c�.�=�R%��}Q$�}/���{�)��#v��H~ڔ{9�a�p��d�L}JY��{5�bi��*)l*���Ws[�`� 2	A���nO�1�:S�xX��i~ HT���/����>X0��B�jB�Jr���=�Ԉ�a��e>����OKU��'� D}��p%=��xJ�)��7U/�$�8��&=��i�է5-�pcX��=s�7�Ҡ�b��BP��&E\D,�(�8����q�c����M�/���3vH�)�o�~��w7I��5j����=���[ ��tZˣ�>u�WR����9jS��^RJ�F�	X>�o����T�DNyXN���G}/:`��e��Âw "U �Zmyʑ@���V�ӊ�4�.��P̽��Dtz��ְ���uR�6��:����+yK�?h�ހ�?���1���h�C_��*�DG=�-���Q�g��ă�-���$���t8�Pى?����tI2��M�4[�2���__����e�I<�/W;uֳV��YE���q���ɺd���9�k��F�ԘK������|��HIʅZ4�ۺ����n��wU;�T5,�d�c�<
��H�p�y����ko�/�o�u(����C�z�bwK�+�d