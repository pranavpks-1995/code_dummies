�i�\7�>������I�$�}�)b0>#V��3a�#׷�w�`<�����8���^��m��e���Q� ��e/���z���e�EZVn|U���	�]���_�S��U�G]�*3��]fc�ȵ�Z
�7��n���~	�'Ԉ�d�b́�&f��r�F!��n���M�;�{��Jc�*��./pK��`�����s�Dg�V@tx�[���y%��j?����T���!�<?����GI�6���[Z�a��!�D:rurભ�>������S�飆�̞��f��z�n���@�R{����/ٛaXj��Tt/d�52�z��s&J�;�.c@0���w3��g; �z�b7_;��4�ȹn!>�}ʞ��]��R`_(�G��`$HA�T�R2Hh�ꢒ��ǩc�	/0�F�)�,����C/�f  ' �F���,t`��"#��3�ȑU��]D��V/�<M�E/���o�{!$��i��oY����������EȤq9�6����2��<�&�h��'=��O����O��_�(���Akr�~��HA =e���*������Nn��];�$˷�]ʦ�F���E�r(����֨	;�X .��m���fNS�2�^~��k���Z���A*I������j��T�f��`��N�<�.�j��Ck;+����J�.���͌uB	<rg�o-�n��;@bd��ǎ����`�F���̆��6
�,,��rɑ�����u~a�
�:�/+�cM{�_:% 
�.��Rm�%��L����c��w�0uAr��-��&��p�$l$��hY5�~#j��Ï��s��[)0|`��4p�]RtT30��W�a��}?�22z!O���[~T��כ������U����ޱ�'�mg�R<Y%�.!e���3#)��lb*n�q��Ql��Pu�#H'y� ��=@W�c�v���	"�_e��I���Cs�n'(Lq�9RTGF��ᰡ���RK>R]6îh��aل��d��氏�H�z%�fK�SOy-ܕ +	�%����%@Uw˲��ZMnp�.�
���x�7�G�2�d�k�I��[�HP f��e�У[���W���l|����,�kO#Y[,���y���?�Fۧ+�d9�8?}~�9�����"j�l�L�.ᙏ3���>��S�9&�G4 �}ѵ|ia�c`=�p� H���R'��SU-���V�`s�P��.���D���   � �-W�����ML���y�r�<�_���am���|@�}O�)8�S�X�,-:���B�g|Q�����1���^�^��ʾ�}���pêqۃK��	̫e��h
��|����^�NV�w\���!P���G}���;mKF�7i��p��X�S>S�.��ÀBA}HѻMy2i�pA�ܳ�̑ˋ=I	0Zƪ�!�к/k����y���U�"��/�iM���q��D�ᖉ(��ٯg<�4�a5����y�jφ��4��@R�c w���[���E�%�Q��_��Q��zw��Z�o��~���	&v��2I/�S+K��"�������v��_͕5�d;�+�Ҳ�Y�oI����{_cWL�y���{��e�Y@\���e��j�x����*�!�h�i� �Js���$D���J���l�$6�זa���K�0�=C�L��u�!t2nM�lٌy��dxG?�+=*w,M�L#��V�K�k���2[����\�B(k��a�!:�F�L��!�iZ]@��b~hIu�5�m�AyH�ơ`z�i2c���h �K��tW���U�XA�2ش���0Ǩ�C�&��~|�fYmpm�fص]e�	�r�''�P�@��_��>��/ّ�C=�J����G,������ЗS5�l�+��lD��0��9%�Ա�����3���I5�Q�ȭ�K���j�N3����ǥ"B�Bu{������>�抯���]��\�h���ɷ�%�_�����E�'5H��
DH4l�l���d�U���;��O�ߚ�ODj����v���A�i �_\�$kh{������\�C�0\(㠦ܸQ8��s`[���@g�I���r�d���I���r�Ҥl�ᔓ-����$�@�w��Ҹi�z��������F~�)�"�8����~/���\u���f	����F0�[=Kco�8V^���7C5bqR�9��_�&�{Ɲh�JP��D��+B�[&;9�}4v��P���
�A[�dLy����l��6Ř ߌ�[��~���|ڴ���z�K����F�����?�����*$S���S��� ="@_�/yA�?Yq<�f�]E��-�Or�?�8!��w�g�r��;�#��r�Aw�b ����m��O,�G�3�O��   ���UW�C���/p�ү�9ʝ��d�/�E�x�HtV&9����g�����Ap>�(��q�h����9��E��� bp��d�jD�O@0�ᶦ�W��!�˨��Xl	v{��
��X�̀|%�̎�O��u��'�!�t<e�	(�
~n�+�r���xP�Fn.�֗��bH;�mdgH��x�Wz_�[i �)=7/�Sx��6�����>�g/�ei p �E+N�:��*o�'3�v_�ya�0@xd5r+�>�Gk%����qjl�x���x1��6��>�EZG6ӋW���@���ՋDr����"}%u����x~R�P�H^���]��?��� �eN�{	���)�Ft�Up���Gn�������F�i��3��u7GEa	�NMv]Qʙ�f�L�0d�����ݐ��v+c�m{��7��xU~���dUpp�ܔ��hõ��9��`f��Ю��s󻎾Seh2ҫ�%�� ��jBgx�36�C������^'�Q�0ʖ���h�*��e~��g"����6/h)g��n�!s1\AG(��EK�cj��bnɚ�5�\M�Ԫ��;9�V4�q�B��EX�/
���%.:�8\]�7%(QwP�V2�H��}��A.sE:�lY���i�@���C?���B�h��H�~HyjI��֥+"�<�-���:`џ|��Y��0���j^ʏeh�F�R�,����+GW�G�o��D2��A�_I2�}�����L`@RHp�
��kC�g���i}�ۧ3�/X����9[�Q���a��$3IZ�n�sIf�϶���#��Y�#΄B�uʬ������r=�[^L����X����@��L�G��o�XVB����ߥ�[��,��TY�S�k>��o�� }��tV"1�|�a�"�n�BSŋmѮ�M�'��(3�S�K��!�<Q-��I��X�V�Y�Xdl*wsp��*�ۏ�U�n��$߁3��i��;@�J��oaU��I�[�����f�e4��D��]�GW��R��D��