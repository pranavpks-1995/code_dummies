(�թ����m�2pr&������|9�# 1��_j�(������ғJ@5�9��ޚ��'�D�S��]l�y�+k���+<r^<�Y"YI�Qg&�E#:
S�Q�EytwiG�8�J����i;p����=?9ﵤ�ˇ��$���"b^������-U����	I�R$_�)_�ˮ�e�E]�U�e��$�Bk�00!/R\���m~��F8��/�.�cW�r��x�d�-�]iJ!��$G�m���6Hɶe����֋�מ���S�t�ڶ�qc����b�tB/?��2ነ���AJ�T}4�[6�xq��Ws��o�&*A����&u���S�0Z��K�"�
�>��sg.�܀�D����7�Ic�����a!B`pG-1�,v�Z,�:�Қ�H���B_a�Tj�M'E�Nj��qx�mٔ4V�#���V(��j���7�Z�����Vj5�LP�T� �Y�1��iZ��I���䙉?�x�~���D�br�)����NE��R�	;<G/�|m�t��Af�/�=���ao�`,V�u �_�����(�%����{�Ǵ��f�5Lܐ{��˴d`���)�����g a�I.�����?��<f��ƫ�F�G@>ް�/�jf�m.e���l�%�NQ�bh�Ox�b֛��f�S��y[�ԝ��%��J&�lX#{	�׽���ɫ�e6��Z{�?f�U�І���L6|��IO�b�' �$ql���n��2�[�;�BQ�x���ċ��� nȅ
H������t�Xk��u��O0�Nv���y�W2�N�ǡ�$9�^�*�n�2�{���珸���7�p�]�C�ޫA䆟؁k�6�]��<����F���v�B�s����m��АH�z���Ƽ4��儱�X|���)G\���	@�q�B�7Zt�@6br;J�IhnԲV�����\U�b`��)Q"��޽l"�O	��Rk��$�@���������Ċ#����BKw����hˬ&1S8UL��:K8u��vH;��^ Ƈ\R����>��
"W��tһ;� N�,��(y�8*��K�H��Es���~�Ւ[�%�A�f �Wz��a؀������10֫��������u�{�<�~/��~8^*�ɠWm���n�h��1p(VГ���Je���8�c,�hx�����O+ߞ����|[����b(/���� ���ge%�����)�N̓���f����	�	�@!��el��Eu�o�����ǝ#8.��#��=�Q�G���y������A�LO��8kx�������v&k�d�v| �{�{�}�>�+҄ ���l�5U8���%F���d�I�sx_����NZ��@3ɥH���$���=��F�Wi�k�(��#�s�z�0\`�զLR��,��ٜ���������d�k��C��=1m�S=Թ")Pk�#�<w��Mp�Y�����F�؁�rޜU�d��	ҷ��	��o�؈�*Zi�Z��F�@���=
nq��Z�_	=Ǭ�08	i����t��} �d�jY� ��Q(E�^���