9��煗��6�G��p��t�-e��7�0��+�������!p���H!��K��}(��V�I1��#��*6���E�їJ��̤�_gs}��ͨ�iW�b�79ٓ�zZy��wBoy����_�0�*�=��<l$���ˆ馡�������V<
��;��oH!&b�U~�{�f�pW�{��X-��-��w�����*�Ẳ�ͣ+����@�W�:���~�k�; ��=O�4X�X�T�҄c�JU�&k�ܐY'i@[u�&������{�Fq�0Z8�:r��� ����aZ-+	2K�͊)���kX�	�Z�c��vn~mh�.�;`� I$e$K�;Ȕ�KD�4W�U#/��θ�<�+
�wI*�~ee0�o��~�o7��c Q�\̙t��� g8*�A��w.�
���� �`f�c���@������~�O6\1�筞���<'�� ���sǧd���hϠ�v�*5��o:2�[�ޡmi�@o���l�E]�k&O(��ueX�{�LCx/�=\�l���W.�Ob��h=���N��P�P{�]�^��OEÆ�����������5f����X{_o�5"l��(�:�]���})$>��Y'��j_��(����
��l������a����h�M����,4�8��e�����'�
%�������lI���%I@.�<q�ȗ�8	��_Q��Ϝ!�HV�����R�Ɉ��-\���s�mՕ�=��[���D�N�����i�5�P�[ݲ�/c*���>�� 7���:T�2}�/9�B���	�� F�n8��2��ԛ7�lf�?F��A�.8 ���������ǿ��r���g���3z�4ޘ0x��|�7�V������>@�C^ �		�X���b���)��t3j��i�Gન����EJ�d��}j*j%�dGf�O����*K7h~o'�D�(�_�Ƭ4��7-�:/mV:�O&�ƣ��/����
aF(�Gy�m}���ȩ^eo?��1���`�B��Tq��z����3����l���J�<�f�Yw;�9��7fb2)���'Ҍ�+"��r��s7�_�����eGʫa}*|e6��C@W�#�N�-<�g�̰���LCP݋�M�k��Ң���������xj�8��"<�s����p_�d}<9bh��b�
%J��������#�-���fj7B:���3Y�fH�Y���k#� gs�y�bCM��5#�r�!FO�x#&;�P�p�� �{�d-;+���rA��S��ߪ�֑��
\������E�>�H�}AMF�@3�P����7s,�s�![���=���2�h��k�:L ;o�͠܀��ط�Xe�W�R�(%�9^^h�5�<d�r."���(�CVD�{E-���P&�r���"����k�R�,�Iy�]<op�~ݩ�ur��S$ݝw�����>�����$����.�oK��q���1��X�"2��\.u��/P��E����9��/���r�2��=��z񲊅!�1/��5AӤ�:9�c���K!&�y���@d��Aރ�WR֥X߼��>�*K���v#����'�����g�b=~2틪C8ip�����t��eB>�d�;}��zu�NH�o �b��6Ҧ��U����jJ��:3?x��<�q�����	r���-Y�q����"R" �* 1 �f�C>�":n��O-��������)]��3�΀�/5/�Y�͑
�^�ֻ������|�k�,���&�z�̩���RDGz���I���W}|['���x�`x�|�F��-�f8�rQ[i�\��_��"�%�[��
��Hde�8�	i#_\O��,.���+q���bef�B�j`��h �=�:��z����_��.W��|�@�6��/���-1*(�Q1�Cj�[���p�1�d��A�өG��"���_y��σ}#���(\ G��9�i��<�v�Z�< U�7V�̻��'#������yv�M�Fi�b<s�{Ϙb�I���@#��[,`��/Mt�EbAr4+�:��E"!�?�g�N쵴���L��j�t�	�.�ԃ�PE��B�R �� =~%���"�u�t�0��9�7����x�D��R ,��:x�7�ůޯ�U���}�9��8C�K�Y��4���K�@F�m��po_N"����:�6���&�����d�ܔ�A>���o X�~�1V�>�,�w\�8s�q�zV+��X'�ù`�c�'tţ�������]����@��?�n@�gܢ��L���|g0��د�����S`�Tp`ls�[R(�_/�Dz:n�*����r�F�c��=矿ΑBå΢MC�M�9��֭>s���rM|"$��q@���|O<��{��'PJR�a��P�Zdl������� cƁ��8�@ݻ����8�"������qd1s�>U@2Q��VD��ir��{�&�S�5�Huޯf�J�� ��yN,[���ft$bB�_g{�9e��{�M���GY����ɥ�D�NN�&�҄[�Cjy�p& �ww�d(~�X�fD����1�;1ͩ���"��ͫ��{�%�x�PRw��ף*lʱ���U�
�Nxp�{r��TȈ�����F]��'�H���jۋ�t^�ڒ��W��wͣ�@��䡖)c���Ø醗�7�<�2�����>�IL�A+Ö?�7�ݨh"䒺F��M��0��� ֱ+���j�m~�&۴�e]m�_[�Ĉ�!g?�Ң�W�U��tLzx{��'�9-��#Oc#X������c�%]��T��y��S��}@�?�*��'�+���>��AQ�i�b"�}�r�EN��9҅kv��7 vb���ݩ��d��&F<C�x$�R~��%7��B���	�E��H=.���w,%�s�K�͔�:���gJe�#lX�M��'(���ê��Ϫ�OpvPܕ[��P��4�#�������HZ�Ͷ^!�#�d��qE���oW��0g�8���z0S�/��r���a�"�ut���X)UY�=F]����(%�M ��X�@�<�UX����H��c�(:!����Ჸ ރ��>{�
2.�����.��	�Z�/%A� ͭ-nֱ�-���xJ0s}����AK`'��!:G$ob$��H��t~T��������~|�)�s-���,m�V.�:�I�%b#��Z�����Sl������" t0~@�C��  ��b'R��c�I�2�|�9�H�~ƅ5�U�P��"MZ��'t+�Yd[�>���"�%��ҥ��Z���%ٵ��j�;��J���`��tT�����S�<*,�c�1'�/��O$'([�紣���� �{������y�=����"e[ςu�� �JY��o�Z�����4��s+<1{��v���Q)hɹ'`j�]�Y��w_��$�3��u��kr�w��o�����VY#����j7�vv�������^��N�G׿^A�~b�'f�z�m�|������џ�Q�������JsV������)�ꪮ�*��tg{f����<�<emu��)�vEh��N �,(���hg�f7=RG<xa�"���l�N�Ƀ�#;��%���d�1P90חW$��E���>��>��n�,�
OY�T������2�Κ�v0��؈��pKʴ3O>���481�k#����x�&i�𡄇�T�v�4z�f�2fQ5�g���D�f*R�22�����4�k�jW�J(�t�c.�}^�<)N/ӞK�q0�zZGrK�rxpEЕ�C�u0���@|ЂXD���$7Ū)v���V�4ţ%������j�P�'���?��2��jަn��Pnw��&������2�MQ��Q��KG>�5)��'�z��ֺ
�cz�5�]�V.溇��/�PX�j.䁔 �J2��"���Xa_a=s���`:�M�t¥�(>�SjN�8�����8�-��� ���'�Y͓�8,߳ �IM#��쳾�H�HI���G��B��(&-`�xu�gG��?d����I:ܑ�q��Ǒ!�\7�]�G����g<���i�L#�