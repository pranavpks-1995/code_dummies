���j����|(H�0S���Y��[���i�T����|�d�?������?��M���	��-_C�ȵͫ�$��m��u�<���8Ԁ�F�o�p�2[lh�ؤB��Uk�Kđ��4��s�U�'��+�#�k+b�Rol8V����p��|>�$UWu�E��ez�Ԫ����Kۮ�RoT�`͌�vw�i�Ɋ��G?�j�sJ�qD�BVp�D���w	�ŀ�����m)B��+��YU�$	�q�o�[Y����ǆ[��o��kI�'l�����f5�N;������J��'d@��[��1��S���6 (���H5��&�d�	�%!t cB9��s������\�IڣC�[   � ��-�����d��LN�m*��ܓx�1��\�,ԍ��<��@�m���搭�@5����N�͘��kmT�� ���0�Ĺ���܋h2[�|�E=�.��x���_p�E�i�1�ښ�����e
�CqV��q�s�s �+�af��H�݀�UNl��fXݒ{7&MT���ù����&��4���<=�Ņk��y�Us���q96K$ z��
�	#{Rw�aRSh�"�+ţ?����MY�:�s��I{�B��׶�3�jy��>ggޜ �ʺ�A��'��>f�����L ������]�T�-�u�!�g������_��H����| ����w�~K�} a�xY�9䒛�.��7ظ��b��k)�����2�*��6w���3Y��K�\J��Vn��u?5�ä�j�IUĤ
�T=�/��p �[�1m
;7w�>b��4rt��OY�@���a*y��q�]3Q�@H���KI'\8��,H6O^����l��!U�F�>Δ��CJ%f�8;X����V�T�z�����v6&V���S��v��֒6;�S/t;R*�����|��y��PmO�2Dy�{�$D���1*QX���e��\�`��g�7qߘTp20���zlݻ�I��ϔ �L��fuZ �k��B^��k���L�m���&��m��KD*-lRbJ���"���p�~R�
���l�\��&����n��Z�8l�r��(��Ǭ�ÈF!�u��9��՞o�d�"�tcU��E�õ1Q���DP��4�-��޻�o�;v�/�5I`��Ҩ1�Y��A)����Sx�(�A�j�4e�M!r�ó�rsN�K_(�l�6�t�""2���?$��g��Q��i˳�ZR{��Ѯ����	��1��$ѓ��V��F��Hq�:}�=��-L�q?�Sp����Ú���]��T�������C�������j�=͋j<��`IxK�Ҙ"�A�Z^��ϋ�K5#C�u#7��۝� b��  �  b�*��\��D`�ϋ�:�W�K���֮���C��E$��~W�^	{�:5��M�b?c�h��J��'7�F!(f̛�G_3Ƿ����n���X�d!����̾s�z�P~�dNU������PLM9��poyYn%���N�V��=�-}�ӯk�����?��_b��cwp����`1J����p��c2����9id��B�x0�јR?�sS��l��Y_G�����3��F?�k�J����K�I'������{�g�E ��({㡛�IY��͗�ļ-���*�X3'�9	�S���KHߴp^�F/ItJ*x�(iWF��
x#��w�����v*K�[�R���	��&�(����f��l9�}Lѭ4ヲO�=}̎j �1��7z�ly>�� 2���oݒ}�֖�-���Z1��eTC"����G��B^��$�`������B~=$��cbl=�;�����H����Bٶ�|;�ʃ�u������@w�x�[�r����q��8Y�q��r�իd�W�p�Kv$8�ߢ�U��_X��?�La�!�^�?��+���[[%3�n��&t-����Q��@�#��w���
�6���Y�����?`��wY�%��7_�+
��|"��vW��:��k>��hT�uM�$Aר��qX��24�!45�a;==S��U�~��|�|U�I�b�Z�<�bz<(7��3�T��|_�鿻+x|#=�m��]��zY3m������t�$NHB��Z��!�� ��!߫�\�ў-(݌��8��:�����?zf/3
�6���$緣J�#o���(Ka��X�TxQ�c��5%� �)�?�Y1�t3�x� ��8<Vz�z���X��-�'�M @�A.��������u)3�YfnJU�-)�\��v�U��.Ϣ=Щ�
�R���B^��w,]7�:��x�7�x��oT�R<��D���Q�Y<�[Q$]/v���GM��`_4��x��V���k$�z�����T+q襋��-U��Q.�D���~ɞ@�v�A�a.�㜫�&��߫�mB,z�N����$�v?!G9Ŗ=I H���%�~6��LO�:����>�vt:�Nc����:�3�V�d�eªl6��x�����l��Hv��,3T��S��'qS�г@��X�_��'�]~���v�0���6��=�au�KB���x�CN\q��[���� `H��>��|Y��h������N@ �'8���uc���|�>�]l�%�|��t���Q�d�� ���.h�9��r?�޳A�L4�zť�k�8��/�94��4n[ژ0{.���L�j��ByOU���ln�W�- ߕ�T;Fk�*�hJ����,�}����>����R�Z�c}0�o�RG�5�
s�'otp�K��w'Vm����}��X��A8��6�y��w��%H�bR�?N�r-'��Y�l6�����=kxH�ץ��Z�69�Aû��I�f�D�d���\�����g�c��U�e�͌$Ϸ���%�X���_Əl=��d�����;b"�����\�Mi��6e!t��G�����٨��j��`�b�~1���3_�",�i��s�X��[*:�<>�zI�9��4c���q�2��I�n�mv'S(�����=��\^�꩗���C��p���.wJ�X��!څ�6���@���X�a'jxڹ�Չ%0D_u�j�����H��=�RS��5�����&j�4�\��"^�Ș�S�E���z�y�X������X�kU�5��h�t-�(����su�����T�\�@s�ī�U=j�MrYr��y��uؖ>�<�4wkB���!�H�N�)�qk�:^n��Ў��;��'V�)ʫ6�ʧ���ch��nC�H<�F��B@)+`��ag��u"Y���,��U{ ���V������~�����c
v?y���L��_�y��ɑ�s,�M8e�Kc9c09ܜ���}W �U�l�S�c��fW��/>w�C�S� Z#e���xcg/^M�tN��V	���'�����Yh)�-D�q�����\���HF���M�X��ʹx~|u;yr͔"jҨ����E���E]ԇg��H�����#���#��M��!!��L������g�nZ�!���Nxo)�Sɲ$���+Bv��w^��W�wX-�By��=�9̈�R�TԴ���]S_on�l���J=�?e?�;:���5u����.f<*0����P)��(3��Jv�=H�F����]F��f��9���ц}���*�d����h"��7.��}��Iw�b�ި���S0Q�� �#���)-b_�֣@�y����W����Wd��&�~�:o-q	ʪ�����@�"y/�>���G��j��;aLOtIS��-0\��=?�Վ���O�� �w�j�$����)^�;󽃶��WF����sY���Y���«)&6��ZJ���\a����3��j+����&Y�{�K~�Iˤ����	@�ˤ�(��g^%�.���G�$��vz�iĕ������ѫ�������F_�� ���QIW��Wg�ݑ���WNMXU�`��,7;�+Q67c�͘�A�0��Y+���y�(�7{��t�x��y�	�9m\}�]GZN��A��9Q/e�i��]������&ʹ0�Xw��/�����Oxg.���(4a�U�N��oxO���1����?W���2�(�k�x�e��:���F~�?��M���$k�YV���m�{�%��&X