e���'b��U��0��F�#k+�R[n�U!֝��Zi��N��*��8���B1}�t�u��2$���k4����vGS�hV�����mп�k$���Ps�z�d���i�|���9	���{VL@!�P�#멓�T`�:�̪V���a��L\Ak�Uj�T�P^���-�/I�����d;�3D~Kn�lc��]�[��G~pJ2�����h�����'�u��B!/�N�����(n��<:�_ȑ�H��%qN]�o1<��,�Y�SG����}=*�'��9	��$�;ݔ- �]Y]t���NC�9~e�u9ۖ"~e��됛J)g�mpΚ&<T,�땗����I� ����z�T ��C�mwnJ�ĲY>�| 쩓sd,�D��Ē�/�a%��oO��dr�A�*��]�,/�Q2�e�#5pL�6���ى�B��}��!d�:�:���akU�R��!P�r|F�J��RG���byd�����[��Csnc�ʑH�&���1��VK�ZsJ�n� )Ȭ�qsl��o9����v�н�8f���8���1��y��g8�~�Z7)���Ҟ������4B���e��
Ec���1����DZ&�+-LEi�������Ca�	�dߏ�MJ�d�V�]_%o���>��,@�a�9�"�)=ҭE���-�U�EHhy��,�l�B���#��lY��u5��b4D�b7�y�9�N*��7������=zy�9�G����^��Sj�_I��\z��y�̫�@�q�W^s�8�(�tw�?%�q���o���wl&uK�3/ъe���4���� 'P�[�\?���f_kxW!cgK/��;y��;RĤҶ��5'Z�E�#�?h�T.<��K���3�#e*�r��t�G�pۻC��]�m_>�Ǹ#ɰ��OF�N_�
5XB�����@��x4;W��|I)���E�H��\�l�����z�mV��w���D;�K   3 �b-�����d�&�L������h,�;$��)z�2DQ´G�?0��nKN�ܕ�e�hL�Υ���c;��9.�&�l�4��`�mధ������r$4���E�g��t	9�Ѷ��&�q:�������qg<��3�Re��N�TGk.�3@5��ct���^���%Vi�R�^dTW!�O�-I��
�ؐ���@f�^�PMK<c �h��ۗmN��H�la
[Θ�ZԒЇ/!|�_��Ob�/,p}E��a|�����\�k��Z7�q���B_�P����"��F��?Ū�, K��t��U��m&��!=%1���Vz�7�-m p�Oe�' "ݧe��da��/꜕�*�ٸ�����V�������d��d$���g�n����
���d��I�rW%�<��Mz �����_�F�߉�Cy2�Q�Z|/�2+�e���G�K��	b�F���aN��e��T�Qdݮ�A�k����kit�ٟ��Ux�]���3C���Y��s� ~��F��\����|��RcP����M\�ժL����#Y�=��a�kHSC�}dkg��g�5"���T�F5KJE@�8��Z�E���l$�/��_I.>�a�f�5���yeFC鴚�Z�����֖�UŶ=Q�񫾝핀NH��NY����,�����Us���k.�uvʩ��~qĤ��&�C\!�	ʂ���C^z@+r��sT!n��E ~�;_�K�7��rB����,�t�{gi����_�����cB���� sN0;�D0���|�;C������Q�O'�~���v�шd����9\��yotR�V�u�$�xr�/���GNy�^oTBL��"��P�͞� �@^��9����F�ZѰ�LaD����?�$��N��圫^Zlڽ/o	b(gtA�{A�Ce-��0�J~s�|�*E�4k�z�������8�{\�������F�y(��u�Rn��,x�p�k�Ո�3�Ĝ�r���Ի�=\K�ܲ����e� U�{��s�-S�9;�mĂ��aU9(r�D�,�dvfܣAR����!��9.+�0 [���y�Km�!�Q6��Ը�<�'e���mҤ�(��XQ���*��Q�ly��"�#a(��������w�5�P��k���(mV�� �39���d���F;�fC�����h���]�|4�U����oЎ�UP�j�u����]�nhff_P �!�
A�("��ob��C$=�
�����>���Ѫ9c�0-��9Q[j��n0�%�\t�Q��)2�,�h�+�aN+�$�Q��l� �0Jj��'|�or� -R	�O�dH��lQe�����`�������H�@�H�
C�Ut�������F� 6�f��� �I���   	��0�W_q��*D��֎����L�*쇏G�(>�@�Ʃ��U����f�'ӉC 7_S��f�����Ʊ��!��=�^X�η7pq�����,�Z��
^�j�S�F��M�\���](|���d0�Gh�if��ڲ9���-�`N�i �K��8�ƌ�n=.+k�D�-ŕ�`�����֦��{����8�a�E�%���÷�UD]���`���A�(��]��]��aQ�w�t�|Љ]';
�zꀾ��}sC�QM^Y�CI0�:���B����@dP���b�p������^l�QF��]P�:`O�(���rh{V�6�ME�E��1�+9M��;���J,����>���.u���>��IA�V;w6�$`�eS\'���	G*�e�6�s��K�U���GR*�*oYR��8��ܒ,��y�l��3���?��k����L-��!���%�oW�*i�e3	p�?=���������\��>�~���ob2u�>���s����Xrrg�g����{A�l��!X���hE�wK^�a���S��#�n��J�ZJ���,A ��ɶ�4��nH�9�^���1�����F�p�i@�@I�AQi<�j�����FIW#z�nt�������?��Z�D�c1(���J�	yh�O{E/e���$"�'���Jײ�p�+�� -�>������ٕ7��n���-�L�9PS#E6��f���9.�����~�
`F�X ���hO�ډ���_�_Xb��#BM��6��h��֫O���9W�jw���>D�ў�J�;)�"�����B=Yd�S k4��r0�)u ��q'F(dү�������i��O��F�{���g�DX�����Jkk]��O�d@ւ����Š��k$� (^�.��\��2��^B_�]Jx���ē/5���#�������L���*ø�$ ^.���.���eѽ�]�����)���MU�/�����p%曻/�n0��G��`�4Y�df;�p�*�
3�� f�6iA���_k��8��JU�ٺfU+���ԑ��v�404͇��ǹ���5n��M����g%�9[�"+�޳
��1��f�@,h�*�
.�z�,5�Q��j6�~�OU���T��RW\f͕@�c�c���	p�,q�}�j��Q���w�F�?��U��ߩ��G�����a�la�'}��$׷i� ��u_