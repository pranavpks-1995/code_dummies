u\('�;���f�0�𔕇��J�>�~����L��i
�ξ�8�c�t�Of7P��h�	d8�2  �_'��@�i��M#�	�Æ��    !K7O��1Fc�"V�8��t�>__�����Ҵ��W]�3��T�[�	��g��}r�Q���5�%z�l�����}���Е�e ��ahqXBQ�R$aԐ��e�n0׼�gK��jW[�z��;BI'ww����{���H1��!��]tp�Zt�4Ƿ���'�M~��     p�K΁B   ��X����C��0!��S�n�jy^��z�:��Z2��i��bz%z��Tk:c�C����k��\9�Fi)�������pVޜ]J��0��E��-��)}Lt s��b�.�\�_�*�s�_��0|̙0+Ȥ��gT`�0�Ԁ�ک��k��el�݆Ω��޿�ѯ�Z���	[�>�����8��<dH���2��Ęx.�Y�T���]�x�#� ���Y��oII�'wu���d�*���9�9?'��&�8[�J'*�D����s�v
+�,X!<�>E�Z�'�π�6"�|IF.ޙ7v���l.���o8�x���u����&c(A�\W��\�A�������rH(Pf9�u�tq�#Xt��A"H]Ad��
����8���}a���m�����!��w+2�Q��x�N����}�"]��.�,3P��',�]����������^��W����y!!'���|���Сnl���C���D��#���(�����Eޤy�o�E���N�D7��ա k��8tk�̤K}*�����*�ր�ӡ�5��)���CGA~���2�um�;��/��#�![�_�N*�9�M��"������X�:/^�?��r*F�^�����l�"��	����2RՒq��]1�cN�����HҬ/�6�1�c�h%Ĝ�w�k]^�u$%z�g~~X ,T2�Y�v�}#֮��T�����ّ��[>��������Q���c��W����чk��u� *%�2Q����	�7�r<�5e)h�}I�\��Z���=�v|���U�e���4�����j��	�Q\��O��:býE_�����
�]����u���V��\��C�*����EK}Ds$+lQ s�����R.��ag��>� ���#q^ ~�BC�-вZ�M�<�!k( L��r�_��v��ۑ7���/�0ԅ�z[B>���]�����19l�"�����
�2ˀ�M2�=>n���wm��]� ��o3:Lp[7ld��Ӫ���ÌĹB�;��H�� �S�%_�'e�" a'�;�zY�*�Ĺ�,�Ĉ0���5�[�\�A)je�'�O�֢�aq&0$�lL�\S�@��a�݅�J�3��w�O�MiS��Ё*v������_g6��Kz�*�i�l��=cB0�>?�Vq�*>a��X]M}���W���H�%�,(u���ks�HѬ&�8��>���IVdYo��N����Is�M�V�̋/��?���h�����~�Q)��o_��N-���hcDdW�6Թ�q�1xp�J�K4���L"���z�qB����B�ÁA˗?M��RY»��jwܻ2
(_�nfx�T�������L�}fhR�֕*D�g���-� ����N���l5��| $
��P���M�t�5C�7����W�4&K�%���,�����o�a��H�^7���Uxlѥ=��,�[{1M�cY�@��Y?B���3�k���JR�VL�tr��GA`-����ކ��v��`�K-�yȬ�1�@>y�% �>h���l� %��&i8��MAGm�̹��qhRt��j3>N���Ň��c�j!���H�>,ݦ�����������4����љ~�/W��mnS�H�P�`W��n:5�CP4Sj4A�-���|��i\-Go�&��o&�����C�?+7:����$<�~�܄��7y<^����>2Y��X/�'��:A�֣�F"߾�fN��*��|#�<����g�yF��p=�P� )�/����F0K�؜��e��[�W����a�}�&�����;����`��ǵ��