;�{��
q7��GM�̳%$'a6�*�.��!����
*spH���Z������JN��j�
�R�"���Z� 2�h�f��d���Z�� **c�&ʝÕ%6�q��A����^a�d$��QB)ȹ��-���U�*�b��I�O������6v|⒥  ܡ����Ӷ-n�α�Izc>�9�����䐏�MM?y����e�nYl��o����MO�Q�ӂ�X���Ʋf}�A��[��˹u�%(lKjY�A'�"����p?�lxI�N�"!��@!"1�(���8W �l��rFwoT����=E���f�m��9m���B�p�,��\(,�j������'���{�4���bŁ�e�:�m�_�F��X���֡DW���R:&WP>�x)*δ  �T�L����ݴ�F�1(pT��Y�O��K�4�;Mǧ�A}>4H��6���5)%-�3���u]�E(z\s�dt�s���D@ݑ�SK8;��<�XH����y��ct��2�
'W�?|В����@� �2���(d�7ʭ���.拳�PI�H �e���s`�M�~8�g��uJU�C��A*0e: �]��1��	��;tu�Zl�'��A�њnh�E3o(lb���N�"'���H�� ��2K��|�����YLz���V��� \�EC�f�5���M�{_�>���׺���_hC^+��z슂��s��bˡ�r���U��F�
�`��U�X+�*���9��t-s��ֱ��~��o��qs��e�Ϯ{�*�C�P�F8��
��*ñx9.L��+�q��y�0��H�ޢ֊�d��F�0ݚ�w	�=�a�]b� �4L�����:�����@��������@�������	����-wa<n�,`��{9ӖV��w� �|Wf��6#~��~&@�����\���v��b!�x�R1�t[v���(�]>���i2��