i��_1��:-�kV?7�U-x���!���o�U37(4���p��0����I~>Km��u�͕4��K
���wN�������@��^�v�b{:2�yxe��#��'��m&���<��{^5�!�R�|&��0X\�F�����ޓ�q���]��;" c����N;�hv)��،�Y&w��#yͧ�!P�Ȕ�1��x�OپgWa�Z�˓u��*�.���|�t��y�N~dv�B�X<�-�3bX���z��<8��жK���BB[s�Xօ����Y����%�{����{��/q@3��a�A���\����`��8�ce������y$S�C��<%��׆��_��mp	6_,�/���=�loV���I�5)hl�9[��!<�y<�J�KZj���Mf�/
q0�5;��#��E�((v�S�=�2޳:]5@�4{	��׶�����8�E��/L+R�7����/+�B+˞�m�ym��{2�(Vč'�u��h�y��鉞`w�h��Gr���>.q��8����v{��Sj���t���}�K�Gh���Yos��k�$ 'X����*�	w��E-���㒄) E���/�︨��S�*��[�O��Y���_{
�>%$HX��P�{�`�Ŏ��+Eo�p|�Č�*���|�H�n�S �j-�h���u��`�VAϮ���+��:���2����.Xc=d�dC(�J��%�&�#�èx[��4�#mb��y�lmq��O>W{Mi�\����{��l#2�����j?j��?ܜ:���wuQ�!/�-�^U@.�?	�	D@?@�v��\K��3������nWv�.OF$iPː��P�߈��^��@��<A�j���(l�,��f�4?��Lu���������.7q+(A�(��ʹ$>�*� ݒ�h*S��lBH�¸w\Bo��=5b�P$�Ǝ����-j���`UGy������M}��GB��3�h���}ru�1(�~�{��uR��)�/�o2�9�����'�3��Oc�yf�126�A4tQ��)U�&�}�;%�����s��)���ֈN.t���A�㱸��\��������1S�G{�Iu�db������g�˂�7������;�m��\,wD�'4D{8�j�u�ZvL΢eG�Q��B�U�R�,D�����a�0(�Ȉ�B���!eH�7���!Wnz�j<�F��A>��C�t!R�$��ݯ}L��\�3�A����+E5��l��ܻ^7h<mZ���mB��n~�K��r�|a�r7���#�6��'��c��h�h��TE�R�8��"�Ȕ�=��}��D�ɪ-�M�/;ė�ޛR�߾�]�����2>�����;'��ZO��3j2Y�5��֩�d��q^�7�j���r�٦�����dF��t˥^;�9�C^� � v^91A�u�/4"�딥�?w�N�岻\/z{@���Y�����R}eHD�L���W�4!o���[���	�D*~
`�+�M¡i�5��sL
�@�Ͽ�r�ž+����$U
�0+aZ�P0�3�]:�#���l*e�F9�r�L�s�Y�<c�Jjy1�W�!�m�;�j�����Vl�K�^�ם9(N�m������Q~դ%�1#;�Ŏ-�)QH�����+h'� �&��l7Y�%?��.�
���r8�
p��x!�e��V���}X\�V�#nƪwXU_���J�ѩ�J:'���b�rR�=�',L@是��;�Ҿ���v��=��%�!U4��h]AlU���hiSR�cd�@�Sě|G�n�󳃷�N3�\�x|�@+%��aSͬ@����P3uq�N$�ر����������c0( ��:���J����pj v;���(Y�&��K��6���Tiω�[���y/ ܦ1�����%G<(<���;�@�`��:��\'��y��툯�:Ht��P��R�B��pN�N� -"�X��y^�d\��>|ܩ ��f�D�SG��T����7Ǌ��״�XO�K
��ǂu[�<p$�fhMLu��h�'�g���é� �`C��F�G2�CҜ�S?�/����A��0HS�)�1�{�_��jh畸��@�K<�8n�o���ZF�ZZA�*���>#�V�/wʸ�|��=�����R�Q�T�;��Dr:e��Y���Qv𶳴���' ݍ�C��:%���A"c�9�^�5`���rn�E�+B6�[�_נ1GX/g��:��o��,RX��rx��8urr9
*����1(�@�e���=;E�]�,��R�yܿ*�#@,#D1E�&r��t_u ��Mͤ�M�ae�<����T�}��9�z��{��izG�e�¶��8\�%��lTb"�1���dr�~e�)0-�h����.��Ju'�`0����W��,f���P��C���Ȣ�*�$�g0��"d ��z�G5����(K�����72��B��H"Ñ��KH;#R=�+�����v:JpoA�w-�B��PNz�[�����}q��3����U��g!f��W]���8~��'Q���D ��}�����}e������?/�g=��<���`j����do'С�UZ oW�<��an��|f�uO��дJ?_K��3�5h��ےn7`!z>y褛�k}�K�:��s3��4��	��0F�
e��kVh��Ħ,fNV����^Ҽʮ����,d�CL�����������)[&M�B�D���'*0M��C�J��/c��OWZ+���}��M�5���,��w�r{��P'H�\��Nkbsg��oA��JE�`�Y Æ�&*�5�POvϠx���Z���w|V�g�U70)���a���~L���Mۈyu��URx��x���@��ZzxԷ�4�(���@�O�K����U�$6��!`���5i��i8E���̠�8��#����{-�\i?�?���w�[).$F����= x�F�aæ�|��!��S�X@([d�_�]R]�'�H����;�{c#��S�ʺ����0�3�j�t�����h~ۮ�<c���7ΐ��"�7ڟѧR}_�3��E�N 
�}vX�����w�i�5-�xv��a�"��I��o�Q�.6�|�#Rp�
Уz*iv"����2F����U��])J11�}y,�,��0)�Dܓ�1�,�;>/
N��qLk����)���� ։*�b��k���	��^R���JQ�#]�i(B�bIEP�u?o�cD�Qf�U�1��lTCf�n}�����F� D"��eз�����To�3v܅�9x9�2ډ��+X�7칬E	ﯼFk=�de�O�$��p��H���ӎI��ڏ��r�TAN����A���}n?&�<�"�,9W	 �����,l��$/z%��-��e���Cʞ5��܆�`�q�
��Uנ��L�Yc�(��ם�/�9���7��sO�A;�E�@>��\9V+/�fW����G���!�ù�hô�=��� ��$i��@9;se�����c�����WyE}Nq�=.�6�2V<����ʻC
�a�9���o�OL�͙���Y����.��̅0�7,�32�l^����t�w���W���-j����j��ڵ@B�=�W� }�����_y�C./:��0?��\O�pLl:�بq�>2�S0u|E��a%�2�LL������U[׿�63���I���e$�6.�Q�/������G�T��ADk�֣�U* 
}Kq�^<�)���-u*M~���������p�����{~�cOSX������+������Q������PP^�S�<�b��!��㘔X7�aq7��	����_/OV�%�f�9����;�Y�>[�<|PH����*��Â��x��=>�31�RǤ0��,[G����e��[¡h� ���s	ɛO�j�%$���� ��7�8|Dܘ8-���͇�V\{��F���Vklr^��&��;�{���cG����n��Ui�����G�	�'X�`S��0���0�z��r 0�eeU�!ʧ�l��)��Y�^M�>ﾢ��7���0(���Vo���o2�A%����M��Sn�͙D2�?��<�<އN�%�b�(��Q17prԺ��hC\�Ȩ�v����̞5V~ ��a�\�@�pܼ�DsFu5����wN�_�dE]D��hs��D;
�Z(�>V��뒦�GOV��۝Z���H53��v��ƹ��E��h� �ѧ�7�(H�/�p��>'&�n����)���1�M�3���2���m�njS�n=Y$Ƌ��� �S�A�~.$��O�n����jtv�\8��؝��[4v47x3G���;�D	��YTn[�� )��zMLx�� �E;3�>�ր ��g����!�-�{=
*|ȟHh��c�ŏ�t���%g�?Lk���0c�cڛRŞ֗����R�=�L9��-��Fv�V�6<��-��RK@��Z�"�~t�f�%�k7�M6���Op�k�����s�k���#uhM�S2�IJ��#'�N�Mԛ�_���Ej�9�����s��߼r����0�������T���)n�	�ɥ�U�D�n,� #���/����CwNO�v�Rh�nˠO����8��V���^��'���@,�e^�w���!o�n��4����t�g-IT
�=� ��%|*�6��ğ�UZ,dJX�E�Hi8�Wg��u����nc��;ǉ�����?�e�~��Ls�� ^��Tp�'��mz��K�ۇa�E��������@o�'��̄]�����̈́�����WG�SXw)��0u2a������\��_�����#�C�u�Y�%c�~��̏4�����	z9� V�G�˻�����!�cF�W¬ErV'�*��v����#�|�4�gy}{R#��
�_�o�G"\�:�F ن��n���+ t	{Y�e�*U-�H(�����ה2oVe�g���<�P�p��9�&����&{��0�>�s�ពB0�?���\������������������l&�^�/-m͌�f�¾��-l1ힻ��Ҹ�����T6�'��q��ߏ��r%C+�Bb�<	�I�B"h���~ߺM���.#TEK{����*�lH�̞��Gh@Qp��"&�s�E)�[�ُ#e5׽�qx�3�;@-b=++ 2o��|2H-^3T� ��ϬĜ��gB�JǺ̠�uo4�����>m��y2�I�/��c_ �%U�?��KM��O��t�Z{�Y�H�T��$��bH5~DZ���oѥ�>p��@%|�k�V/`��2w����7I�!���ҜV�VVw�^y	I�"�n��JM�o̖��y,׸����\��iB� ��xT�JW�"��~H���sw�qxۀ�N�|>�G����iވ2�[��jDm�Ŧ"�x�㍊M���W���H?bԱt���-
X��꺾/�\�{_����q�%��v���!�4dk	����%�G�~�fpC^�ޙ�;�ۋ��� պ��ݣ�����)[�~ޮA�M[|S�!ׯ��yܼ���t�6c����x:�tD�I�6rV��܉4��������˻�$��pts�����捓�Ra�����E7��ұ"��ܕD6}��8�+���|8��l�ֻ��$�W�aՊ�|���������f8	&�+^IO̍��Ã �	`̾���a� |0��hՂ��� '� ܳƃ�����x"�oX0��H��Y[Dc�[�U`�S�C�ȕ�k+F/[(��T\�O��h���ĥLi����?�����!�(&�/,�Q�����GB+��˔`�MoLbj{iZ��:���m]2�.�>_8s��F�S�}�Q�y"J2��N+�EQSA!{��4��np�ڀ)+;*E]�IVЁ�+BEN����0�����Ȋ�r´]eL1�='1���Y���1��0��3k^2�Қ�Tb����~�f��1Ⱦ��G��;��q�j���]��e<��f����3o�G= �2�w�U!�����-ֵ�&oQ��]���?e�\FH,�n���8��n햺Lly�M��I��h��P�;`����5;�K�8��%�1��$[�"F�Y�Z6����q2u�w����X��Z}'[����Q���X>1���q�8^�����&�m�pPh�25�na�� ��r���|1������J��֫�fZ�_�;!�*��[$r�0Ji�^L��q{XT�^�c�y�2���v%��l[ёU,E	}���|7��K�����|�����E�� �����Ԡ�!��ă�hl3s�F�P��5�]I�]��]�X�!|�����|�n<���d�@�S�mg�rL�Xa��J�Mi�%�R�s�<�=�%��$'�z.o��K"|=d�O��3�t��ie�����f�c�E�x ����! ��Zo�ۧL!q��:B�N�~��{�   !���A��#
n�X�$a� �3Ŧ��u^~"2� �@��x��'�n��ԡ(����}������o4�/�j�i��I� �_�a�.���/I���s�t�*VQ�E�D�8� (/#�0%1!�����%�V�)+�)�ee���!��i�� $`�!($�ۄjtD��l]�U i�H^Rϵ��qD  !��50!P X e��=s��� ��n��nXJ��>q�ʚ�fǫ��"��]�����c��.�X�k2�#���5���S�+�]�|��7d]�=�/0L�e�e�f�	����ee<�X�v.W�ٴ���g*&�t�l K+�2  \Al%�'/���cXI	�7����x.���m���|Y	�r `  @0!)��0�2ţ��[	V�:.�21��]���h��������:�������)���eyZћt�.Ǯ^�R�W�Qک�#� ꧅@�	�� � W��J!l%[ @�����Ϡ�����s�O+%%�"b�:n��{�]�£�S�c�T� 0�B-��Fn����HbN:�0    !K�H��R"�ĥl��A%AXo΍�)��k��נ�ҲQx��1B�)�����-�B����������pz4�V1^q:UN��������������2��ت�-`:X�+���A+
FD��]��Ă"LSH%N�0/of�lA�@�`pȐp��z�����>�K���q�����T�<�!�u�%��n�Q۔�'��Ӡ    �!y��0`�D@�@��   �"��S�㝽Y�H?2qq��O���x,%wD�_�>��"v���X|���Q_���S��aK�JK�+�1Tn1cTѧ���׺g��,�����	��Q� @������@�{py��Q��T�O��t�����     !���6H�hC "��ă���Y����5>S��hG~拇_C�h�m�ZEt8^g[ _������h�"�\�4`)t�=�H��ZS��/	�-��W�cu�qc���hu]m %u��J�d9sΑ� 	-��b���ٯ�7+���     !����5���R�����Yk`������X�ҿV�ؤ�HB�﷦�$�
&�)�BZ�xͱ� ��EI*�^�C��d�84��|R)�i��M��\��(1�j�	�:кU �a�H!�v��b��B>�]#7U	����\��    �����  She guessed 8, 9,
based on his drawings.����J7� �   
/��I�c�ݽJK�ȱ/D�������L��<�7�b�a�<k��1�a�8��2�+m��*�0�uG԰ ���#�Іx?�5]�@�@�+Y)�����8�c9���}�[��ǜ�0N3�� ዽy�00�"�k���*�:X]5(>G�܆�ێ��
QY�6�OO�r�A§��=��҇����m�o��;���Jm�k.-�����$س���WE~}�D��lHƺm��.&��S8�� �<�׫j�.G��$l�w�ݭ܀��rZ-�?!�*h����IP�my)��*�;s|��[�Ղ�L���zx���a�,~ʣI��M��T�2��)�����!
W���{����3�j���t�����=O�J����^��|�q�a�93����>n��Ǡ]^�+C����H��1S�p,�IYČw�n��5���1Sl�����-�lדX_���S�$��g�������d��L�@��l����v�K�����m�+s�uTZ8f��%�+���3!�6]u�I�.a2��y�~r�h���?���h�[O60��/�,�K����ȎX� ��b0��U�L]9;��L<�j��4��;F��B*(f���M��8]Ђ����p��@�J@0}Gҧ,�"�������{�[�dmq�ڢ]��yS�q�L�t���*��֗i��P�6����N!���*���hn~�Ɂ\�Wn���i��C���>�|����uP>aB��W� �����X��H-�+i���$�����i��=����<	��2�z��4��(�%�}�a��?�c�cL�V�(����mY��D��	N�e�b�Z(Q�*8�Ux��ע�J��3��H;�ż��N9 �VJ�c���9�
;[��!��wR?~�y�b�n�zR�\� Wȫ�Wɪ|�<E��r1IT8�v�{1f�3ZvF\
v���k�ފ\"B��{�gg�Oj<���s�!���Y]���EQLV8�aAg0�l�wᐓa��}�z�'�۰����:���s/�ܟ�Q 𒷪�ӎ�~^�i���b!�f�E�i�W�rt�椪.?j�9:��_�EyU`���ݷjG�Qc)���0é������Y���#aBS�@9ƫ�G} J������=������{aM@�E�65�"�Rs<6�-������cu�M�jȷfJU�igj֞/���d�?1�k�
'vFãM��3�Ĕ[����lloc��i��*���t�'���F*�prm7rDMU�vuj���ň���C�q ��� 5���0��#�HQ����k�����g��nx|���p�P�n��X$'d��H���M_�?��@рlB߫o��0��hB�}��fċ2R����h�%��~"�����'N�����Pǰ@�͒)�޷h.��*����9ܜ�Ob�&�0�s��g�� �vy�-��[%��ء�����O�
6�Ĵ[z�����M����Fb�J�;��A���#U�E��:���oa�Z�>��X)p=�*�
&*D�B�b��U�3�G��6��79폇~�F�I��u���Q�J��ږF��윿����ʁ����rM�ҧV��'U/j����!�G�(	��i)'}�;���R@�����������݅�0�Δ��-�z�-C�/Uj�h:TE�)�zI �6��v�r;���O1���ȯދׂO��~k���S|�FeJ~^7@[��\C>��6��b�ڪ
��x�xR�k�H�=;��r#r���|G7&��t�D��.RQ��]w(��ܜ@/%��6�E(5=e�� ���$��C���
�� 'd�V�@B�QwSY|���hX�-��S�5=�e?;RӐ!�p9��B�RǮ=��UX��?5L�c���}q��c�=�g��D���V-%�?Ce�k`������.D'G�-���x�j�����M����5K�p�'�jTQ��	!Jr�nߍ����C]�~	�w�&�9̇}G]h\����=���q��.H��❶X%j�&�_�,�!.����B�⅋��� �T��t��O�,k�݂���j�C*����M6���h�6\���3�ޯ�L��5��9���P�z��'��a����`o���vw��փ3�z:���b��{��2���ic��o5cȒ�̕���)H����-G�:9��*oȖ/K|�$囉��駺_�v�h^��Og��@�O���o�t�O+���;��Z��"�Q�=tOo���EO[_=�J�`�#n�䅌�R^`L�?2�3�����M�G��Aݯqq�7k��4������HԀ3�2����|EО�Q�<��Xw�\i���p�hȬ�0��dJM�?��4��Y���ꇋ�*�H�qr}�q��@
6�P�6@v���[ǥ�,�g@�U�:�|����@��w��]�g���]���	��[2ƃ�K�+AHu��0��.���ͲY�<ٍ�} �ʱ��z�&��������j��ae���-�����C�� T  ��xc�wc��ë���@=d/���0C��ہ�wsI�ܒ�7������R~��Slqonx7Y���d������Qc���Ob0T���th�|<z?YY��9X���W1����7�s�u�S��MJ�z��@�+61w��#�!sR�<���{R8���%�v��_��+�.-�0��ͭ���ت���K��3.�D,ec��2{)�+xS�v��CC�u�-kpk�祕�0���D��������f�^�FC���#���}^?�s4����ؤ�7GYz���Zo�9�Y�e�梮&a�����0�U�Q�}���$�%��> �����֧��Aм�[S��ݍ( ��c���Y�r�nAd��VrC/6nQ��W�N����1~��%Z��ۼ9�p؀i~|������ ���C�2���M&����P������'�x��J�$.7F�W�bi�����)�uw�:ƥ^�{}M`s��5�'��i˴|ZV��K�J��ٴ�I(����y�o�E,�v�5D���R��U�4���W�ý~��M�!`g؈qEնr����.� ze�i)�&lk��5�o���T�f.vpE��8�'Q��酂�!��(=� ������g̅���歚s��!��f�OQ+!LK�R��ו�����B��pkm^|.Jv�uR��kݬ�*���8�ߤ�N���H���T\��C#�ȑ�u���C�];#.#LA�'*k��@��T��J�/�=#�`u�Еo�L�@��J�'��zf$lb�/s��Ѥ��d��B���P��unG#Kk� q��78�s}dU��P�����:�@N_CΤ��0-o��g��U�N������]�����|&�(�B�ܤ_�}�`OԆ��KHCZ��b� ���f%�t�\�{�j����y�J�@������12���toDS���}8�\Cn�+�Av�nE��nW���6��_�i�n�{����g��9
 �|W)O�s�RI���.�A{� *  s ��~�|/��,hh��C@ē�l2�(%�7Bq�T���TA��߃�q��8��P�+�4��#��r_�}���ji�]-%L^f���l�b0���qT8�i���Tៀ {mx��w�`�`�\/5�� 8 � Lnpj�;�8L���'3�xG�,O.$�^l��OhS��S`��+t��6���G
�+, ���?�����$yo`����� �IZ�W�8(�B�<ɜu�]�:u�G �vJ��g��%�@T�g1c���!~�
�؀���x- g�@\�L�cC��W�{��P�և�j�08N����l��
q`vR��>^r�E8��Xy	�b�qw�� �jA���l��` u-E� )��sM�9&`�B� ~    �Ƶ�F:0Dc�� �hhHH4��|N���FjJ`�L	���Uz��b�/p��qWD��C
�^U%!�/�R���Q���*�:�7��#Y���jM�kF�"1��'Fvc�A���Ժ^BS�nYY�u�:��RL��*�J5���*B��E���f��f"` uv�"u�}�ةږt�?6��<�EE�ܟ�_gpm���@3�2��H�N�^n屺��_Ƈ4k��zEr�"�#^W`6&���8�������?yAz���r;̠R�^�����"3��� ��%����z��d_�A�)����i���L!]�]ZB�n��?	7p>�WV�ݿN�����*�C��J�@�ߊ_~��ݶ�g�?Vln� ���5�M;w�0v�w����0ۋ�������e3�:P4����RAߑ+l3nؠs�k'�z�DBc����1����KF�o$�ǡ�%R�D|�o�>��?�tA��:��~Z�8dW$/Ȼ}�sX�E��W��������!��������* |���P��j�������+=��P��~v}����	���*8����J�Q�n`�2�N��#�2�����Nq�'�Ү�4���n�F�DTH��vڦg��|-eEA1���!a�B�y�頖B�',U��X�T򻡐P�Wa��<D�Ѭ��V<x�n�����O  �!�����"0Ц�S�d2�P J|rj�ra���kg8���� D�$w�]t ��ۄ�I ��i?��TJ����S�.�?�W��������S%`&�Կ�G-���e�����z��ޕ��9ѷ|�@ Ҩ��m�ˎ@'DA�x~�Ԓ몢wM~�k���v��U�@     0!����Ac�VEZ�4���+�,dË5�F32�����5/�Q�ӽ�m:J#���ڸ��0.�e�v�pE�����;)@Lk������su�~B��6�����+�c(�1������>P'V�]4��M��o)���    !��8b�`��@e#�@v�r�d��d�A`�$��'�<��-�������DH�:��C�Q�#+�ګ㞅���������ף��e'�������;ַ�����F�g����'.1����;U.S�
�"���d�A_���M��f*����w����/�m>{���L;�]�  !��4�kC A C[��� ���.:m�"����k���bG;�� 0�z����_�r����T@�H�j�(��t���W4�ȁ�W�&��(���鿕����5��0��UEO	��X>��49 �$��UU%��:�V�w�Ez���UqP�;w%� !)��4��! � �6^a+#�I�)�`l(F���^��H�︄z�p�=,��XX{ m���Xڒ�t/��O�:N�a.�J�0�B4��db�V�f�@�=��^5uT�s�
ɚ�J��� �l%dr@�ח�x�����7�i�1UM.�Q�]�H�  � p!K�GBN	R,�Kv&�8�Q� JPr��,�Yb�M4M~y7�\8��h{�����\B��|x�� �,e����@i�����Pk�$�b�>��ي`�� ���Tܩ�9ײ���oB�:�W��Bh*��XTG��޴q���W�ٚ�QK"����,㏘�f�2��ckl@����{?�$��TX>˦q;�`�jO٤ �`�mDP �!KmL-J6�ad�U&��b
L��Q�Pe�'^��(qv˅ep�³ b�}�&�[�9�(^�b�����2�cl��JF��/�b�L��QĹ%˒����^��4�6�z����~9���:2��=z�u�N�@{��X ���4Ѫ�`��' �����k,Ul�T�j�˅   �M��x   �� ��}�0��M�8í4{��5@[A�LH�׏���(���s���42��S����Ї�aE�;Nɧ�W�{"&�*����EڮST�Zr��ۥ@�� ���h��sn.�:6�$Ӯ/c0���7���AB��y%h�y��ᄔυ��1"� ��@�D$�w�A0y�S�p�*R	�ڢ�+:��x���Ȳ�9����(ƓKB��@tG|pN�����U��&�sp}Ymq�83�ȈS��.'e"DS[�_�ɦ�s��H�j��,P�FB��Bc&Gqi� �d����m��F���\Rت,�e���Ҫ�R��3
g���$��V?.����ރ,o�o�(%�T_g�)��)qȭ�m����d�]D@��e��߮#}�:Z-zVp�>���Q@�w�1!����n���W��c]�yl�3�Z<U�]�qj]�\�y���Q��M[�'VT�!�8��i�]Z�k���6ce��2�Кo�T���"�6xJ˫�W� u�v�-~��%�}��L��!4� K�5�SۡI�,�_�&��2��UV�C�h�-H;я#տ1w����j�ֳ�B������`zdT�m�Il���q6'��H�Xs 0��X��~�����Ò�%������en)�lBZ������'q�BY�3�b�'�/��F��T\.t��b�ʄ��G�^up�_��OC�4v��2XQW�K�.*���D��Aq�`g���_�� �֎��h+�w�B��n���R:i���[��'f��0:���G,�ï�������' -�}Gk*�d#kx�:�7G��f������Ah���c��;�N%�e�~�t��k�<%���>����'��~i��N���vfQD�Q�5�:|�,
T��� �*�S���u�dV*����� �P�ή�*��%�Y��m�MM�U����X�ş�\nE��)¶0�<&�-s��� ��?^@;�g�WBx��(��@�[���G �.�Cթ���PP%�FVqK����T�,���v���\ZM�
����>Y*zՅ���X�O�l{�L�|��$B �I��Bam�[�)Y,p8AR��^���!��0:��q�l��N��eL�
z��
�g�����8i~цd����y�<ݛpz��G[,�{b
k w����;�?�b[V$&l�Ŧ��0���W�|N����T�Z]N�������QRS��
K&�bSϏ��"J���Γ��6Ũ�m�1Cs��� �L��&a���`|4_1H�~g�l��8�@).�O�~�]��Q�\}��}��T�� |��_��2��}��I��Xy�772���x�0O,{1�:;��\��l$��J�t��$��]|�BJ�ľ��V����7�[ܣ�w��8Y�{%E$����I�"�")"�d����̫-��ږ����0���a��M�cq7��-��P��>k⥔�h� cƓE��Y	���c+�6�_��"�ǒ�ź�uΦ���g��rN��1@h�?#�>� �i�y�(g����t���I����mH8��FS���6�u��/���O��xr7yL��2@{������zX����S��;�����*���[��l�e%zós��ٛ�w�o�p�6U=���Mh�/Q̐8^��j�_,ZX0o+[��)!�OX� j��)	�Ӿ�PC@�����#�l�M5[�&u�V�R��^�	�qh_tH�ޖ�(��R��;oXW#JI>��\��9'_B�n�ߊdW�Sc��;�i��Ƌ�L�^ �8'T�5
]�肿W�N��J>yD�����d$�kQv?5�ڏ�m<?B��z�)��#�m��U���=EEv��cq��e��}�eWd�#j�(�1�y��p�,�؏�f����!�E�y�ӯ����bhN<�Xs}����%�)��Y����_��#�
�T�n��S+��*��_(�:�U=�J�H�¨�Rx1�93��[���B-e�EY"s Z���SX?a�I"�)'NB?������3I�J%M����Ŷ.2>!�kS7�l֢P��/O��nL�Ā?��L�\�t-�)�;�:q(�r||��<���$��8��̭�Q�v�������m��ݷ��cU�@��~ɚ�I��wfF��z�u��^k�_g+Q�c�.��ABՅ��3i�8hW��0��J�-�:���DM��ܺH����	N�e�̏��J�9ޣt��I�!�Kr��E��΋�yޛ�����UۚhQ�V�@R
����q�W�)_�=[l�nV躡/k�;������2^���t$���1rf]�bQ�o�H��%v3^b.CV'��2�[*��i���`�T9i��I�h�)S�-ӧ,�� Z���oR'Y�bz�I��(��ve�v�~hD�?����|X���Q�	����cÐ�b֧KW��[�<w�����U�J���ȧ����q������SS�A:@򕎙O�5����V��q���Ys��<�qջ�~,d��g�w����X^`A�#�ٹ4�̃V�.���C���/��NM;�7H��"������M�nλR/!��TP�M)P���*�1��dI�c�=ߞv_�����3ƌI�HSp��c8_���ɼ6A��qŖ��|�����i��������̣.��߳����;�MU�
�����T��q�@���`2�{vI�1�Щq8a!��$��m�[~��m���պy����G��l?+�9N�a�í�
��I�G�-�|�X��MԀ��PB����l3�+�C�k�Ţ�m��c��.��2��Jܢ���7�*��Xb����o�<�.��K�7��R^��ls��sF
����QL��OV̲�������ζ�ٱ���&���=y���x��u����r�l*���9j`���
����9Y �"��[�h�49�P-�L�9�� �;���mV��;���#Fp�}��ٯ�8�=|�T�+@�%���ZՍZf��t�JV��T�.�nx:?wʪ��4�eM���ab��~��y�)ͨ�fD�dfCKF���&�V_:`�x���Op�n�q;^vM�~}E(��e��4�&�ʤ^�0��$P�KD��LK�4�BM��9��h�X�ñ�1`Q[��(���KS0q�ch��I(����fP�{K��C������D(9ӗ�p"6��L�Fj <T}o~؈�y8��@N���{���lOB���Q�̖0���9��t��&�O(�n��gW1���M%Zder���=���`�%ӘN�Ɉ�hB��_�\̑C烝��,ێ������c<:#�D��t�+�:-�K]'ι����o��O�����^�L����G��6��@�w�5��=�8�WSʠ}�D����׾��Q�n����E>��'n�ה�CN�$  F�B'U_q��Z�� �26$�.q�2�����h���@WQ�ήesZ;*�6ʎѽ�:�{�:�����h�Cd75Nm��F�$ ��{�d�zȭ��/����K[KJP/�l�EO%ċ�ꅾeRU��s��;�S�gݗm��1�쀻�G�u]({��i�2Z�[�0�j�т�XĆ�/P.H�&��'�S���05HE@㨆�4���0�(8]�-�8�\�X�HkmN��>qu��0�x�{�{
5��|r��mF#[��hY�?@A��c��Jɇ���(y��U�H&t��3)SrI)_��lv���5j�nL�|��fU�S��;o�~�iS:,���Tʠ�Fd�~��?㾝��R"1!%c�5�5�R+m}r'��x�k��`��L��'5V���2��6��������f֭��8t�9a Q��/o\�FB�n��n1��8~e��	����Ö�kڅR�8�?_�Dd1���.PH�jy�U�,�p��.,�jH(ul��chT��{#���xEi��9D�����艟x+�P�m������[ ƛv�W[�Ӄ�Ѕ�l�$M�S��!�p �Vҋ�Z&�?�! W��mp�c�o�[E�'�C�C�!��k�;�����^y<3o<tԵ�
�a3�P��s��j��:��!�h5�H�dL�.R¶�O;�T�;pWZ�͍�8m5�O}��
���	�Ł�G/MF!#n;�FF`����CCeG1Q=�*Wj�2 �>f�o"O�_�V�z�\���X��آ�XFl����~�\���U��d^�c�;K��E  XX��j�YL�O�Bi� �  a ��U��W.������@�.M���ֶ��t���g7�+�ep�I
�4��>�����2{f�Ѝ�W��0����#�:J1Ŝ�