(y-��$����>��1���c�}/3�����g^!����� I�iGAi��dV��6m"�1WR�X7FX༺(孨����/6˩�b�9������׶:�-0���L�ؘ�}'�f�� �'B���-kE|��|�rh���yku�U������8>��6�X1 ��YI�f�K�N9�E<�v�v�܉U��~�RlV�;�CGq����{l<8ڦɡ��ƿ�Z�@�ቷ=.==,O�G}�UX���?�ȟ}�M[0���b����Q���~�b������ޛ,ŔZ�+��;Ԇ�$�����`�Ca�@~���	�KD�;�O�R:�Rc�!��I�䏳]Ah���H�����5�R�U�������'��'?Qr��L��-����_w�ď^e�:��Q|�d�$.I�kFs�u>��F�f���zYv�0|1\�&�U�E��y��R�Ac�E*r��=��[�DA&�T,���r�X?�޲>���Vo��R��t,��خ��ɺ}����|��~�sQ,��mAѨ ���^z\^��p�΅ۚ6��M��i vy��k��dv����w�Ę�/;DZ��P�g��\e��՗1�'/�$��m̞L�Y�\���Ό�n�l����a/,�k5���q�^Ƃ+c�6`<�����z�X�4Iffo8�9f��g#4`T|�})l0ptTu݉�ͪ�͝�P�BV����ϲi}��BŔ�e�>���R$��R��%��d-'ݟ��jo��������	)V{�N-w_����cbMa�g�NI���sdD6�KpFFȌ����M��: ��H�n��������W����{F�_�5z� g�r�r������W�/D|�8��)��2�#�ˏ�I�jǴ� ���R��i֫^�cϑ{��D�I��eT�k�h޴�j�d�ݧs�Ņ��W�]�B|2+]�y�E|�4Å\�e;���lC��ĉ��(���� �h�U�^���g6������r{���')S�ᐔe�#�����{�O�[(�u��bz���@�52��#j��X���� t��^C���&\�:��d�v��ar���E���p�ṔpP��E��\A��4Qׄ�-��v�FiB�I�r:n�'��+��˴�<mZz!���{�mhg�m�S(vF�����L�"�P�%�_�2�G%Ǌ��V����4{1D���8*� e�f��=�(�b<�~���p�KJ�$��gc�}��h.z�a���K*��t�~?�Ca��9��*����Ac�t�˘IA����� �-Ƕ�p�j��>Q�t�W{����}Y����ئ��c_����ޛ�̲�H酻�`b9Āꃒ�m���C�>�)2 ��%���n^]���{����I�� &��o��]�Y���R6�I�#Ă��OQ|r��=j70�b���pE���41b��~��e
�!�b�P�CP��FơТ �@��s��6�����0t�`�I������I�+%4;K�{�x�V0�(���x������
S������*.�9��l�Fdfz�q5�����*�\
�F����ꏕ��ߌxr���S�d�\򛈔i�V�7^�C��L�xD	z
�R�,�s��]�>C�)@������BBcfW찞��Α�{�Q�$�[k=�u���3�Fx�%��߁PƠ���Bo��Ҭf�I��R��1i������������$A��b�*�?��_����B���vH!��<���b�Q�I��r���]^������ס6�q�SyJ�'�Rކ˘wp��ȷ� ����R�,^y��M0=s���Y������S���G��>�}��2V����i����m�Bm��Q�jva@s����_�H,��	>27=���x�	��!ϼ_gf�2/?�gn�c�;���i�!�oWw;�֯��にv$J�Hƀ�i���n����+_! ����Q.r�@(z�\$�#D�{,�hz�Jq8㮕����-����(�o������ܷ]('�<cg�U�e|���z\7[��	c��Ϫ}�9��)Ɲ�tʐ����Q�^@�e���
P��y'F�h����>��J� ϯ�'C>E������;�a��a�z�z��	�����w[[��"7/U��(j��ѳ��g�4�U6�V���Xʘ9��F0�dY7=�A���1|�f��@�����J!~a-*�8��C)�v(E4�$����ۚ�[<�~��-�H�{��W] Y��w��S�=&��Z�?�1�-���v w�JXSck�8�v�S����=~S�l��g����H�7-�lg �ġ��^��4A}����Ҩ�9p� I�UG6�P�pɻ�vJa�JT�x=��Ѿȋ�5EM����;j���M���p?����kv2��#*!,�?���%HTS��LgPoVXg�M�N���.ݴ_�B�����)����˪,��dz�+�<Q|L��<	;�w~y0����dB$�0��P�al�kq�%B�;x�@V?X�=����"�+�0��&o��髪�v�~��g�«����v�U<�t'�K����k����~S�&�r2��Դ�CD���ъ�%�j��J�>�@�
Cc�7h�=�=�-��g�hnF�/��$�=��9�͜tq�˪x�D�[�-K�Ep@a[�>�^|� :Ɏ@�Q���s���W��>:�Xl��)����Hd`Cr�ߊ@�2���,�"�ʗ�1�:��	b���듧k�/|�|>v�
^��-��o9ޏ��_�~��>Ur/_��~h�(��逡7���Afj���|!B�H���iMm�ZbT2��]�п��ߓ�=�|x;{s��϶G�����żYx*)ϾYčx�x���'D	ќ��me$lo�hK^�P����Q�O[J�-#:�,T�)m��@��hM��#��c�M���\q[���%���ʥ¯�V�O�Ch�x,��X�&˺i���`�UJ�ݜ����j���ݓ��0�ӏ`�9�9m�-�{�c���2��Uz��4۴H��m��	y���0Q����"����)���}j*
M%��3>�A5�i����Tx"���W5͡4��������ļ��Ӈ��^��1����M"G�<�8y|����~�c��s[<,��/�;����k�{�,��;�2�����W*q��XH}Y�(5'�j�5)��+5l|����@ޫ��@d�"�B�n{��<y_�z��T��Uoٻ<4R���J��x)8ɣ��8�r�WA/����b�óF=$�V�� ݲ9��;�?Q���S�+Q�-��I��D\b^*.�����BGz��e/ܪK�����[��8�����É��b�T�Z&��q�� y��^D�i��p�)�d�u�<�^��֌�=�"l�P���S����oQ��D�$N8��Fem��@��Q�9�潬,r���1��a"��P��L�t���=��(Q��=`�c�'\�p�{�����9ì�:WV>�Iӣ=wd�R�D��1���>����V:�oi�J�U�i�SM���А`;	�޹}B�烆�8�t�I��B���&�쁾&In��585��6�������!��#�5�Di��KZ�n�D��3�}0ַzx�5+�(����R�E�W��Q6���_���@�B����&-���[�X�ͅ�D}論8�7���#y�33�n����Ag��p�c�\��$�CS����ߨ����K�J)��O6�V���I��.��]#�y��9�M]�v�͜��oq0_`ߜ��-�E1_�xn��&Qz|����}�"U��4��[���i^��}�U	�3���-ZGH�c%\6�\�/�X
�%`�5�Z�܏"5�\��4RO��x��� ��o���!��[�ˁ���ϲ~.��LV&�1�g5�:���E�!�M�8?�`U�KR��E�a���-�*Uo�fG��H#9����,h<^�����-u�F���Qm
]q��|}^��~����	8�gX}|��I��,�+��u����
��f��7�iC���M��7�p�%10<�:�D��UE>��:L\����l���+r+Gr2�8�� ��"�Г�����K��M� Y��K����`1?uټ&�k���M�aгk��N��
�0&�P�� Ug\x>rɛ㣉�rQ|zlW�/���z�؀�7����O{p�}�Ih�n��+�T�@Q��A1'֝�y�
����~ܻ��̋�}Y����b]y�}fr���ĻT��y5N�����?�G(�RE���]8l�Қ.vY�얩��o�ٜ�����`����!.�.��,.q�.�3�(�;G�j֒��w�r�ǌ�g��t\�{{���ץ����^L �;_��cR�i
��/� BҺV�M�\4�>v�2UG�j��Y��N�������d�NsFAoQ�&��k��J�h��{�Z��]��Q��I��! �m�ñ�YI�y59o�1�����Yճa��m� �L�G��l���=��;��O��:�>�����S�:*ъ�M��y"�!����h"!�k��I:�Ė�M>R������t`�s:#%��POXH`|4Sz�~�Oy�b	���P��<�Ş�ٰ�e������I���k(���?��a�^d��:!�su2��%h���r�����/�/�0��o��b1k�s4�t%���>(��o���+�b%�(�����Qi�s[`z'�]|��N5��f4����P�c��4Ꞩ0�:��|q���x���{�_���8d�_�d��� n�iJ��]��m�R
>�!�PLc殩n���j;D��j!M=�w��#�R5���r+"+>������:Aʬ��[ho:7�=������<Ʈh���:?S�k���N2����ʩ�!Z&��,.1�]���N�R����{BR�e��t2� ��G�|��d?	���k���}�8���6��� )��%�ӟꅱ�Vۼ�P����y���1�ٛk,��L)�ѯ�:{�b��h��I#zRݖT��)4��ˬ��9I��]��x���$�����c�Ѻl4S�Y�H7���}������g �Q=;7�$�>�^�t~�8�t���Pj����}Q5��o�P��� B/���KHoE��%��nZ��ܫ�-�ȫsg&�R��,�� �=��#�TĞ���'ɥ�^CE�1�,�߅�IE����7���*�*��|x�%�7�T��~�L5R���Dl�~���:$6,L\�Gc� T  [�"'RW�c��˧r���;u�I���9��I#A���:�>�h ���V�~�S����l��$��^P��<V���s�?���V���M�ȩ�f쩃�=��G/�+8�*3���"v�5B�u�ٯ���dm}k�Y���@,�H�k.lN�zpT��'�0�����!bt�����6���$�7�O�,o���A�N�y'���HW�8�}@V/��S��9O��b@�Ɵ����Rqd	�B��)��8B8�����,���L[�;𛻄[}]���-'ت�6n?k��Er=B[�-� �S���'�G��^���N6N+����
����5��`����*��9��U��٨¾�%��5]���وJ�K�	p:�\��{�F���#L�ъ]G���M�ﯚ�+7fE��>#�&ޱh�*�/p�*���C�S'>�����:5kP[�Ș�:iZ�IPV�aC��EG�'��@�����s�ӱ-#�� �k��XkZ>��5���ٺ� p��:ץoS�gDj�s��S�����+��_ D����Va
�!����Ay/3^��wK8��nǾ�@2,�4��G26~S��4c�4?P+MKR�������P�G(tk{K�A��W��O�!t�q��90�]D�fb�#���<`���	Y|��Y���8)������KU�s-����� �vL~x�L0�?�q�fg��D[<&y�#Uk��P�6(|}у]�w_�t�����3!���!a��CB:�#�g��T�|j�7�>;��I�dm@9�M���.�RM�:W�7o�x.��c�c�
0_��Q�>�}��v�����yն�EJq &����K|`wo6ѣ3uϰ�*N.�(.�;&�e<7��x� ye�9��;�Z<{N��y������O7�
���j~����q:�<����_����*t�(�!��G<�L�U�K�
Ո�=}=j޵��
��0��������+�����؜m F��&���3�:Y4q@= ��m^�K����*�EL�;��J5	j�� 5��S��sj	}wS��:��+�k�M`�4$�e�$�jK��ϣ ~͹�I�	cu��h�f���t�@FFd�2|��n���������^~�g�}��R��Ā����,|%Җi6��c*ç���@�+�w*�./}�D�ͬ�3v�{o^��Ұ�Ɣ4�l��e�J�]�����_��[��+�g��"��G��H���jy�w�������PQ{����i<9OF85����s�������=�Y�?C��:�:%̀�~��t�����\<*��ԩ-�
�0�?�߃�G�8Z�� ���q�}�ϓI�0h��6���j��C.�.��/����P�����͙lg;��u+�-L@l>�d�t^�J��$޳�{�Q�2> x�m���2�cVk9���o�[�K=|[���ݰ+-�*�x|�/�W
�D��F��È�)w�=����Ӣb�4S�MC�y+���4}����~�Br��g��F��-cqÎ0�;/�'}x�+9��������Z�Q�Q��kzlm������D��c�AA�k^����I[�Ļ*v&a��'�o�WOPm�aNî��X�z�	�:3ǩ���5�|<�/@fp!1k�,r^�f<��c�yէ�~֑0H} ԚB��ܣ]��g&���@��Z,�T�Iڿ��<2���]qJ�RE1uW��d�x:-��)����:t`Q��f�M?)��5ר�w�� d�]��=n��7U�0��]��7�9W{��)���@\��@�d���^�B��Pm�B3��^&:�Wˋ,Әa�����S�B�qL|%uˏ0���D�    ����U� �Q�!"�-��R�;$�K�:p0I��X�h�������ݝ鰓�c�����+x��[e��@����n��/�}#/b1j��/ڀ!���Hk=J�\Wʢ6$+�l��)�";�pa�ה�ve� ��ț��K�I�2�7w�c���{��I���@ �!�Tr3XT������.-���3J�����aNDx���`������İf.8q��\Wt�9�#�*�gyn��*��.]Au]�dw��%]��:�a�'�����k�}����UrX�wn�X��wx�J�����.�2����'N�Qݢu�M��55=`���i�G����D�cF����^��l�q�F;�:'U�k8�oO�TO;��0�p�_���W�B�̨!��v��Of�S��報��<즗�����9)ǝ3�u��1���$��_�«�G7e�gg�:�iw�'(��n��M�f^��'E�^޼�c'st�$�aiY6z����S��t22kDM�I_��9�s�~+�A�BrD5��J���xYn���T��{\�GY/�_�'�qK������K�{�{l2�97�{�A�(x�F{@��t�Aj*���)'����R��@�Α\=�F�$E�� �	+�7�s���_]��1qI��a2�^/�2(S���^w�
%W>|���C2��n�%AJ�+��f׼A}3=�xeK0�Mߤʃؗtcg��ރ�ݭ�թ��-���[���w�e�q�Y�t	�5>��V� ����=.wlÝ��M:X�`��x�`y�_(J� z�o�_�D{5H.�qmL�Y��r��ǚ�v&�^p�O5D���z��Rݦ{�/�o���VyO �6B��r+�0�L�d�qH��U��2|9M�,X�Lc��y}� �����c��u~�]��w5!a��Uq��1�4y:rh������*���'����"�FcikU8�D��};�E@�Es�y���y'�