�ES4F�	���i^F/�{�BS��YK���*c�I!1��#��D�C+8rzʷTɬ���5�gLi��2dމ)�¹�j�>�hCY,y���#�fPݓ�T�lG�"Z������h�0��k�>��Y��	���̜>�6	��)D����S�߂OGP�~6Z/&��?E��z�%�T�Y���������k�J��1�g���`fh��VPfH&z��G2�X�@���"d��WX�K�9H�s��IG��9^�UN�X2W�0��C���Rr��Qٖ]5��<0���Sv4i��?Bؚ7���w�F�V��&�ؒF����83���'
�b�B&� ���k�呷:��%6��y�Y��p��;BFyN�L4H�˘mk�<�Ҟz'F-P��B�b���D�z�+�9����ؑ��?�;�]7$��	I��뱘☤�6��a�Y`�h��}�u4��5¶��c��o/*�T	p�U�Q���B���3~�tW-�dԨe�B�x(���v��P ى�J�S�I��X��ː��;t��P7��4�ʠ�xm�#J��Cf�7��e>�C�ƋS�x;O*`�^�"r1�����2D��JC����G
;�5���W&H�׻�%������31<��\�ɘ.w�(.R��++L^磈�<�����n���-�*�
"�w����6��i��s�~����y���n�d+���Lƅ^1
���s��9Xן��}����
D���Z�����	$����B��U