\�o��eud6���zc8%N�Q�K�*֗H����IS�G�@@�Pd�q.H3���K1����TX��8��2 �6N��3�ޝ�K�7\�BV���Q��l��A}�|�M�u������,�KYw$CcSYb���S���z�)s��x�����Α���Z��(
/�����2R?�١���Q�`�3�Y:V�nJ�y���뮁��	�ejT�J�A<�7�Z��ᮁ
1�(��9U�\a��[}ɦ�!ʇ��y�����^8�%JE��l�E�"���:�P<�j�0xwe6UEQv��\lԩ� t��M���1R�Q8�����A#7����7|:���xH�����&��
}b�15��t����q~��&��Rg���U��0�Y�G7��z���;̾���(׸6K��=��m6�J�8��M���3�y���(��k��z��b�����uiU�K�
�i�9J�R�FL4~Ё�bp���ܻ~;�udР��fE���/9�C�|�����}��QxO!�>vlCW��鞃��E�Go�ui�4�+�
���=��s$�#7���s>GpBI��~����A>�,lv��ѕU�T�݆ʛ���(3�.��Ka�VE��4�ڰ��w\x�mヌ�\-7ˋ�׀�"�]gfh";��a��],8\���n�MIС�J^���JS�LN{A����z�;�t<�=�Q���O��)�$˽�op�8b޲Ă����� �C�hC��e8 ��*x�m+�PR��^�����l��5��6�X2����9]nF���E����,����V����*TE���\��غQ�yB�}=���]��/X�Z������g�B~9�}Ge���[�>��}��I�V�'a����kmT:��*Q}#�<���9wF���v{b�[-��4t�B���Y��Y�w�
Y�U/�u����Y���V]���㈷�0�ŉ����?�jCRet�?��ު%+�]Y	�N�Q��EN��28(��+�C��h�?�6��f�huގY��V�sⷳH|1��Q�A�hGp�}
Kup�#���t씶p�!�,�&	~*:iI53��+d�	G���\ΟyE@�b�{��IV�K��ъ�Ǉ���h6R��4w7���!Y��jn�B�O��I�� ח����q����N����e:�6��Aq86 �W�}��-I$?"±���i���M�ҧ�e!u���j�Kܱ���yWR�<�)�Y�@�,�x!D;�1?����J?3�@����D���>ȅ�K��)68�ʊlߦѺ�
I$Q���/�)OF|`y�Yl�����<�4�;F�i���֛Wz5�Z� ��$��\�Q��!���R.!V��ur�Ƌ贝�z�.��]X1lT���U`�I�����X��%줠�ĳ�����uoKh
��U_��=-(�/뚴,�dzJ�_aզOnk��޸�`�z��!PC]�͵N\�՟�v�����p�O<%I,B� ������_�.�~
؋1,;��c���C�~� �E��a`�f=�%Ϣ����~E+�^��}d=�|=�0�M��}p�m�Ԩ"	�����Q��� {�;�qE��<Աi�Ka�;5���-��DX{a$5��k�e��8��]ȽY��B��R}�d�u�_:=W\���~��z���v�mec�#����1p�������ߟj�Hw ��w$$�;r �qyl����ܾ��ΰ]����M�'(x�mx�(��B�	lU➽����9�z��~����t���?kA���V�������o( �g���P��"�u�fy�"��h�#g��A�+֚G�;���l������$��v+����0$���M�x�41�"6�Ƶ�<�J�2H#g�IU����C�T�#-�QI�]�����t�ջNC�{��.΃N��=x�[�����n�svz�����ODUW�;�	�ܹ�
?`��yYd�����e,fN��[g�����{m6˵����A�P����xO���g����-˿a~M1�zU�g.N!���i5�"e[9��5��~�&+�Y_X���x<���uG��*�7�5����\�j�* 	L#���~m%����M�u��P*Qiؘ���?{�����8�?����i�#��j�W�+�+daڃ,D��*��B�bupR�I�E��ge+P��Iu�l���{��3�_*����Ҩ������s"��/�ȦP���f�2,zwR�Q�{&�"T=����6Ȃ1�u<~ɝ04�N�����;]XRR����১~�'�U�sw��l' �$[�fK8{�:�������mih�n�%�+��n2/e��B���
�	d�r�Aw*������BDrs�B�')`������35/�y��Yަ��K��5��}�$?���ш� ���Z�M�M������$pص�x�~4?ٝI��z���0����}��B�Ew�l�U
��^6|��ʣW�	�^�Vw�Y"Mg"e'�
���55�߼	}�5y�@p���c�g�yE��@&p���$�c�����߄i��6n|k���X"������8��a"Jㅜ�[��\��/����=���F�L�
Mj���bHy|*c�xMf��g�i�MKh#�����^���8�[y}����m��r�����=�((�Yr����v�S��G�<�ݚ���}�H��
�B�֥��߫g��ta�R˳7q�B��\��ߥ�d�$/�� �i�֣w���3�R�%�����[��[�"F�P2�{����(�lp��o4'W�6V���=�d��Rqo(+�򹪽'���r�Д7���I�n��=�5ʚ��@��^ef='v2[i����5�5�wvq8�±��7����'�g�������F�T��M