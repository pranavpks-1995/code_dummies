uiaUUB}z�r5班n��^�9���e,R���S#�i��g��?`�{�������n�^5���E�my��m��4GQ�Ũ�~z�9��Ј�8'D�s��K�F~�#�����&��aԂ�	w��,���� ����`z��;J
>���_��JL]dP "?�� C�l�Z�9Y��VPkZ3�%�,}f��gp@�̓Cu��&��4��o�o�Ʉ�J)�p��0��>m�3��9�"�s�Ko��ӋR0_.4eG�4��xT�B:8����g/����;�������$��ϫ=+Ϡ����
ت���\���{�������b-�OG���C�{x���j�vHg�;��xȚ�o���C�/���U_�U�����<�%�� 	��S�]�If)�5&"ۅ_�@ۏ����|�v��
l�P5��>�Km�LI�[q3�rU���"5���Bac!Α�L���<�����֝�?�H��j������9ň�
g��ܫTody= $A[�	�3���T��ڦď&��U��sސ�Н�vV�}�w�#�q�K�1�A�蘱�ɢ�L�����h�SQbWX�L]�#�ev46��%����&��y��p��gq�q\`���&��#j�#xry�9���{`�~��X�2�1��,~�p�)z�,��u�/[�y���}�����۠�G;�*�»��h̜�%��60ֲ1��3Z������b�����BR�ޘ����%}���1"d�@w%�44,;���㑋�>1��Pg��:	Z@����-ב��;�*�8n:��oE���Ey?�:gͦUdk �{/��kB�#0z�W7����`.�;[�T�ݪ�hf�� �ۏ�
��k��{DGm����R�Ҵ�p��M`W���H��^����oF��&
8|��T7�O���;X����@����fh `�+��R��N��|Vr%��%�9۷k��yGUk�	�e��^�}_O>�1���v�N;��k�ܴ����*����
w���3<�M�*a�͗@q�g��q�DME�8����t�u�会9L��O)U�j����)0ߌ9]�W3g�Yǟ�=��¼�N*(b7�(�^�g��