�t-@H�A���~c�� 6)Ǥ1�#&�]�ެ!��%���?QU�>IS7��d������kK�mb�k�
�$޲ȝ)ŅI�� g�6S��*Cx;�{�
�]�_�<K���� �����q?-��������*Tv����%3�Kk����K�RP�1�C�4U�-?V�DE){����A\a�P�oqk����^|Q݄�4���v��W�'@K���e���:�arU�5w�ڇ��p+���ƶ+S���<U
��*�?C�XD1�(a7
�pT�i��Ĭ� Q�3~1�o�|V�ܪ֒J���Q����-g�8���V�Gf�͔� xky�2�J�cw�;��Ť�tn O	�n��ׁi�8ʗ��φu�z=&��k�g�y�>��9S���+�m�Ŝfc�a�_p��6�2S�iܣ��gK���uņ��?B�im.7�,�8�f�^��G�{/ǐwt�7�ܙy���Q��\��ؽ��F�)���GQPꠃ%)�6�@��jmwa�w2��l�9�{�3υ��I��6���@�l8%O<ħǐ~ ��x���6���BS�Z���S4�����ā'����6������ţ\��G^&�����fp^Y���yI���T5.-����V��s�1���&�'WT���A7�k  /�b%R��c����K�&X�����%ʒos����3I���! )�
e]jI��k�\�ɿ�6�Z�+c�h���Ȉ���}`�(i%|s���h���4uW�PwL�txL6�.5kr��f���I|I;�vn,i��Լ �М��ao���.��Y� �@�	$� +{c��6�(��βô�JE�h�u���K� wr���OI��+%���	������zU\1��A3A��2����V7և�G��J`tA�v��܍�y���@�j.we�+/�L��2k��\�S�b������'�c�����@B   � �F���,ta�<��8a� ��!OAxZW�v.�E�p�/�xz"AE�`�����x_mhp�8���r�,�s9)~#� G�'/S`z�����P�B	-�_�aܠF�(n~	��b�A�6��}��#�h���ls���`A��frqf�jK��v�^
]��ғ��蜅�����d��`���y�p�@��    � ��-W���P�F���$p����iF'�l�+in��1!��u{T�C��%�Q�n��ꭇ�8%<0�f�GY�@j1�����
 ۚhu��i D���'�z��c���-k�*$���A�6�4m�]��/M�i�Y�jW�9�+��>b����+��o��t9z�o��-�#3�+�ZˀU$����y.sMb��6~{ څ�=� &��1�)v1�_��A��!���!y����B�B0ozn����h>]���D���o^�`Pi�N� ����b[�T�!�ZmX�vu{��Ϸ*v�-����-��9򲠓��*��F����_δ/)M�z`~� n�O�č���:ZL����߻�%w�r�� 0   0 !)��HaF�*)���aB�x� 	��귬�������=��}��挢����O_znR���'󰇜URW�(���D��1�B�k��^�V0�pE�޷��^��=��� �GM�����-L N��aB�x� 	�����i���ꛫzó{xEt� `       p!K�IBD�u"JGR.�� �m��[+/C�ZdM���J-oM.V6k)�<�F�/;��5|)7�n1�j�N6d����� >Y�v<�[訊�N��_���F�+��u|0�U����B���'���ġ	Tv�}�;�XrvdP�a��Hv�F(�|#�M���g�U��p�V�� `    �D��f   ��ȲUW�D:0G\�{�"i�yT���Ƿ�{��^R�5d̑)Н L�(�5�̓+]11mY�ʹ@����L�	�â	g�xd�8]L�
���^H1ri��w�h1|��x)���os��#����f�{QL���\co��lj�p�.a4VDboz̔�z�˻�ⰑCA��g�'�NFǎ��ɒ�F��-& Wa=,Q�	}��]�jw�#�4���/��(�]=g�mV�zu�ש�l� "
gS���ꖬ�	�X���uע�:{؊�R<}��*s�B�c�Ĕ�R}�:L�]a*R�3���ހLv��kѣL�z�zt�$�M7���-<Cgg�\�s*@�=��I����l��y�b�l����L*����p˪,h�ȴ��F�9G�Ȑ���:o��ך֤d�ӝ�L���V����,WL�{I �������ZlÉ|��ן}%�2E�o �
\y���j�&2R�(�`Q�{Ҭ��@V���♪u���x �j�����ڐ�Ñ@��̀��e�f�a��Q������\{:�V���%�63>qK_�c�3��$-��4f�nc��\绡�۹��<P�A�6���瀂�7 `6��a|����� JD�#��hn� ��R3"���C�r_�[:��Ļk^�|�Ǘ�<p�o�u�6� ���z�تq`V"c�f�����0E��J�fj�u[\�����������, �n����İI����JYFE@\�5��65N�en�x�_�%π܇���6�.�&fO̘'��ҋ�s"Ǥ�ޟ�#��-�R1/�c�y��JN�8kT��9�d�^S��z�S1�#a�^��� ��[И�I�~��|%<t�pN2^�mw�|)�1O�?�`.�_|�W�S��?9~�H��]�Ouȳ�k\�z�t� �я��3��S�'4D�bѶqB���{�(�ҧ��%8l�%{���.̓���qL|���U�Hs=�76!��l�<��=�8-թ]_�>7��:T��)T��Z�c��F�h�v#៿��Љ��9�*<@ 0Ϭ�v�X��b&Н��%�����
 ���& ϲȠ�F<�a�Q2���3�,�9�*&�-bV+]U�]A�t�k�`r&��ۙ�⢭	|��	�w�v��Á  ���%RW�c�	b���'TP��P�U�3kj�b?��������t0<_,�B�A>I\�og��u��`"����:�#}�@,�5��M�.;�7��"�A�%�[�Z?��(v4�t���^�Ip_w� ��C^�W�z��	���'��:�{ޫ:�Q9�o��E��������	�C�����\<����	��I<�bU�R\@���X~(��i[��`��|ң�*�1U�E���1�
���B+6ˉ`�ښ��7W |ؔי�p%��<�đ?�>� �ޔ���W Vn��ϔw�]��{p��YC��@��x�%$�:�E�*ԯ�Ȏ�+;wi6�e��:��