H�H�x����6�����B/�nS�=����A!8c����cI@�(-U�tM�܇t�G�p�z>n�>ED@�ٓ�1!�-�] �Kr��ǻ=��՚����?T�hӒ��c\I؄@�1	͝�B\Ve�p��Rؠ��r���&�a�G�DI���t� <|�9���~�q�$�u�� ��	<��=>�� H:��U����7�#^N��q�d|D�>��R-����㋇m��b¯)��W����J
A4�;��H_�\�b+A�o���޳5�Y��aD��2\3��C��8��򫑾������I��؏�{�Eɲj��v��8��0[�v��G��ѳ1g �5K�}ԗ��j'D����FzBl����5\.N�/���$�?���
TB�Q^,o_be[E��]�un��No�v�*#{ ���6����I[�i���v�h'�}�4�E��V��jvrl�s������R�Z2�<MF@��D�����DE'�Ba�g�N�$g��L��ӈo���p�oe�@L��6���~siExO}��B( K�4=dԨϏ+g�
h�T�ݼ�q6�I�\�t��m6/���.�FЩ����he�|L�/TRp2�
\s�&��o��c|�*��h|���Sǰ�n���9��6h��U�XG��`�� �;�����\�d�r\ �j�[}��l$# �Ф�sq��)����t��!g֙Xy�)�`������Uh򎶡_WI�%��u0��B��w�pB�ڨX`V���ӊv5U���+qj�|�Bp0�<�OF��_���H��h7�$o��L�o"	�[�OM,S:Oc�����~�Z#/}˶�)�iȒ-����(�݋g���g�� 0�V�u���Dk6H�Rkf�����'��(TI����^��.�U6�3���J�:K�yMN��z��IfCd��D�y5?in���1��Փ�g����Y��w�#V��|��[2 �'�[PwJ;S�1�;��q�����6�&���:C�Dm;�x�-����>؍*c�ࠫ�L�����C�,���$���]\)�?������0�z�@��_j���`�H��	�   � �F�u�$4#�KFm�f���m�N1V�8H�]��> ��HH�g�e�ZV�_��,���A��K���)<V��Fm�P`U2�!���5{A[B��<"�.�����O��)_]7gi�e��`a�Q�H��!�O�H�e���o���*�`��Ā���������ݻ��R&�ۘ쿦t�f>;�8-�]�}���6d�lk}�W*��?�ۧw��&ɞ��^�ʂ%*��;�4aq�ժhq`c�)�����\;Ί���"��]{�~�����,I�lذ/ϸ�x"��ۇ��c��	<5��?�e�UȌ҄�d��S>2e�$���x�'�C+o�����ə���a{�3V��� ��Q�(
�l�G��Q6�}� l��b��Μ�%.�|��I�zWY�c�^�s��FttT����`�2��cWݞU�K���{��������@?�Z�T�E�����'�8_�w@����Nk4��p���񣩵�b�C��������/�GO6W��S#d�/Xp�Dck_�ϲ��|ᷓ�}lt�_�K|bkݽx�waŞk��_Y��(Y/վ�0�Y}Uc�bFuy-�>����k#��?Qp�-aX{�f���1W�'�zw����P#�2�a���&��^�T٧��x]�[��%U�;pD�X',�g ����M��/i�xj�)	�,�r�N�pz�F�e��/)X;�
 ��Q�H��= st�I=�F$�5�^J���)N�L��3�N����W��=l_�n�2�+uh�T	��+ݔ�.S	N��q]6�x�	�ԏ�1��^��/O�K?�	����/���,Ld�v8��U�2 �Z��LipY��!9�!r��$է���O�d����w ��|�H.J�(1������E8_��z$��R'�'.�ɜ�֤�eV���ul}Duu~��H¡C�zI�t^�=�G�k��S�Y��{�*FK�T���a��}���
WK�Q�O���~gnע=n���u���eI_az���O�LM���""(7rE�� ��a�°�>�x���h����#+�U2D�3M�d'���)���o��<[WSX��j�3�q6�hmd�R�ح��> w$c��l��8��O)�Pn����D1�h��=���$4�L
�g����:yg��o�D��B(D�Z��^M�'+�B�{q,Óm]XW��3�wɍ�ʊٱ?Qd��%�3A:�5ɫ��^�}��j���͞�����s� �r���`���VI��AnΉ�#�mN���������VTOߓy(���Mg�����b����i�Rczgn���>����,~>���]L������s���fɼ\721�1��.�H��MK��0_������;�=p�pɱ��F�{��j�Ԡ=d��V�S�(�+a֘���!i�`�Օ�7���%S�A@h��=�V�b����c���Oar�I��y�t���?�!34�Q#0�IWE�A�<Jd�+R�f�K�'�
��9:ů�������M��FV��#�E_��N՘8����]��[}�o�j��+Gp�
)��4b�
>�)A�є��9�K�bi _o���n�8R��g����y��G�k�(�
���z��<P,៸'��h�\�=��ИbW#�Tn &�1挥��zL��&�z�J���	Jb��4Z�B�yJs9,���B\bK��5���lm�\��[>����@��t�A�9�Ǳ���L�~�_E����S�S�/�+*�LE��E���i��dZ7@I��e�7eQ�kbG5�(�1SxT�]�ٙ�r�V�"<m������[��Rǩ���][/$2�Rb֖B&����8�,п?0��&p�xE2ة�J[G��#w��իH0um��
Q��gi<BP�?�8��,�r